* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lcesd1_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT lcesd2_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_shield PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_wos PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT rnod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_x_40k PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_x_40k PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_x_40k PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nr36 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_w40 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ICV_72
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_71
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_70
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT padbox
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pad_out VDD DataOut pad VSS
** N=25 EP=4 IP=1 FDC=96
M0 VSS VDD 7 VSS N L=3.5e-07 W=9e-06 $X=5700 $Y=147100 $D=0
M1 8 7 VSS VSS N L=3.5e-07 W=9e-06 $X=8100 $Y=147100 $D=0
M2 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=13200 $Y=147100 $D=0
M3 10 DataOut VSS VSS N L=3.5e-07 W=9e-06 $X=15600 $Y=147100 $D=0
M4 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=191300 $D=0
M5 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=196210 $D=0
M6 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=197780 $D=0
M7 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=202690 $D=0
M8 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=204260 $D=0
M9 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=209170 $D=0
M10 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=210740 $D=0
M11 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=215650 $D=0
M12 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=217220 $D=0
M13 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=222130 $D=0
M14 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=18000 $Y=147100 $D=0
M15 10 DataOut VSS VSS N L=3.5e-07 W=9e-06 $X=20400 $Y=147100 $D=0
M16 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=22800 $Y=147100 $D=0
M17 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=25200 $Y=147100 $D=0
M18 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=27600 $Y=147100 $D=0
M19 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=30000 $Y=147100 $D=0
M20 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=32400 $Y=147100 $D=0
M21 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=34800 $Y=147100 $D=0
M22 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=37200 $Y=147100 $D=0
M23 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=39600 $Y=147100 $D=0
M24 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=42000 $Y=147100 $D=0
M25 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=44400 $Y=147100 $D=0
M26 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=191300 $D=0
M27 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=196210 $D=0
M28 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=197780 $D=0
M29 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=202690 $D=0
M30 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=204260 $D=0
M31 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=209170 $D=0
M32 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=210740 $D=0
M33 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=215650 $D=0
M34 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=217220 $D=0
M35 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=222130 $D=0
M36 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=59400 $Y=146950 $D=0
M37 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=61800 $Y=146950 $D=0
M38 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=64200 $Y=146950 $D=0
M39 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=66600 $Y=146950 $D=0
M40 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=69000 $Y=146950 $D=0
M41 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=71400 $Y=146950 $D=0
M42 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=73800 $Y=146950 $D=0
M43 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=76200 $Y=146950 $D=0
M44 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=78600 $Y=146950 $D=0
M45 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=81000 $Y=146950 $D=0
M46 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=83400 $Y=146950 $D=0
M47 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=85800 $Y=146950 $D=0
M48 VDD VDD 7 VDD P L=3.5e-07 W=1.56e-05 $X=5700 $Y=165550 $D=16
M49 8 7 VDD VDD P L=3.5e-07 W=1.56e-05 $X=8100 $Y=165550 $D=16
M50 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=13200 $Y=165550 $D=16
M51 9 DataOut VDD VDD P L=3.5e-07 W=1.56e-05 $X=15600 $Y=165550 $D=16
M52 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=97085 $D=16
M53 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=101995 $D=16
M54 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=103565 $D=16
M55 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=108475 $D=16
M56 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=110045 $D=16
M57 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=114955 $D=16
M58 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=116525 $D=16
M59 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=121435 $D=16
M60 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=123005 $D=16
M61 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=127915 $D=16
M62 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=18000 $Y=165550 $D=16
M63 9 DataOut VDD VDD P L=3.5e-07 W=1.56e-05 $X=20400 $Y=165550 $D=16
M64 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=22800 $Y=165550 $D=16
M65 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=25200 $Y=165550 $D=16
M66 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=27600 $Y=165550 $D=16
M67 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=30000 $Y=165550 $D=16
M68 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=32400 $Y=165550 $D=16
M69 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=34800 $Y=165550 $D=16
M70 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=37200 $Y=165550 $D=16
M71 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=39600 $Y=165550 $D=16
M72 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=42000 $Y=165550 $D=16
M73 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=44400 $Y=165550 $D=16
M74 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=97085 $D=16
M75 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=101995 $D=16
M76 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=103565 $D=16
M77 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=108475 $D=16
M78 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=110045 $D=16
M79 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=114955 $D=16
M80 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=116525 $D=16
M81 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=121435 $D=16
M82 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=123005 $D=16
M83 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=127915 $D=16
M84 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=59400 $Y=165550 $D=16
M85 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=61800 $Y=165550 $D=16
M86 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=64200 $Y=165550 $D=16
M87 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=66600 $Y=165550 $D=16
M88 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=69000 $Y=165550 $D=16
M89 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=71400 $Y=165550 $D=16
M90 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=73800 $Y=165550 $D=16
M91 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=76200 $Y=165550 $D=16
M92 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=78600 $Y=165550 $D=16
M93 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=81000 $Y=165550 $D=16
M94 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=83400 $Y=165550 $D=16
M95 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=85800 $Y=165550 $D=16
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4
** N=6 EP=4 IP=6 FDC=96
X0 2 3 4 1 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_69
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_68
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pad_in VSS pad VDD DataIn
** N=24 EP=4 IP=1 FDC=96
M0 VSS VSS 7 VSS N L=3.5e-07 W=9e-06 $X=5700 $Y=147100 $D=0
M1 8 7 VSS VSS N L=3.5e-07 W=9e-06 $X=8100 $Y=147100 $D=0
M2 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=13200 $Y=147100 $D=0
M3 10 VSS VSS VSS N L=3.5e-07 W=9e-06 $X=15600 $Y=147100 $D=0
M4 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=191300 $D=0
M5 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=196210 $D=0
M6 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=197780 $D=0
M7 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=202690 $D=0
M8 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=204260 $D=0
M9 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=209170 $D=0
M10 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=210740 $D=0
M11 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=215650 $D=0
M12 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=217220 $D=0
M13 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=222130 $D=0
M14 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=18000 $Y=147100 $D=0
M15 10 VSS VSS VSS N L=3.5e-07 W=9e-06 $X=20400 $Y=147100 $D=0
M16 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=22800 $Y=147100 $D=0
M17 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=25200 $Y=147100 $D=0
M18 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=27600 $Y=147100 $D=0
M19 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=30000 $Y=147100 $D=0
M20 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=32400 $Y=147100 $D=0
M21 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=34800 $Y=147100 $D=0
M22 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=37200 $Y=147100 $D=0
M23 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=39600 $Y=147100 $D=0
M24 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=42000 $Y=147100 $D=0
M25 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=44400 $Y=147100 $D=0
M26 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=191300 $D=0
M27 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=196210 $D=0
M28 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=197780 $D=0
M29 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=202690 $D=0
M30 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=204260 $D=0
M31 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=209170 $D=0
M32 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=210740 $D=0
M33 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=215650 $D=0
M34 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=217220 $D=0
M35 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=222130 $D=0
M36 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=59400 $Y=146950 $D=0
M37 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=61800 $Y=146950 $D=0
M38 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=64200 $Y=146950 $D=0
M39 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=66600 $Y=146950 $D=0
M40 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=69000 $Y=146950 $D=0
M41 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=71400 $Y=146950 $D=0
M42 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=73800 $Y=146950 $D=0
M43 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=76200 $Y=146950 $D=0
M44 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=78600 $Y=146950 $D=0
M45 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=81000 $Y=146950 $D=0
M46 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=83400 $Y=146950 $D=0
M47 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=85800 $Y=146950 $D=0
M48 VDD VSS 7 VDD P L=3.5e-07 W=1.56e-05 $X=5700 $Y=165550 $D=16
M49 8 7 VDD VDD P L=3.5e-07 W=1.56e-05 $X=8100 $Y=165550 $D=16
M50 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=13200 $Y=165550 $D=16
M51 9 VSS VDD VDD P L=3.5e-07 W=1.56e-05 $X=15600 $Y=165550 $D=16
M52 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=97085 $D=16
M53 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=101995 $D=16
M54 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=103565 $D=16
M55 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=108475 $D=16
M56 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=110045 $D=16
M57 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=114955 $D=16
M58 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=116525 $D=16
M59 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=121435 $D=16
M60 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=123005 $D=16
M61 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=127915 $D=16
M62 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=18000 $Y=165550 $D=16
M63 9 VSS VDD VDD P L=3.5e-07 W=1.56e-05 $X=20400 $Y=165550 $D=16
M64 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=22800 $Y=165550 $D=16
M65 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=25200 $Y=165550 $D=16
M66 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=27600 $Y=165550 $D=16
M67 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=30000 $Y=165550 $D=16
M68 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=32400 $Y=165550 $D=16
M69 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=34800 $Y=165550 $D=16
M70 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=37200 $Y=165550 $D=16
M71 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=39600 $Y=165550 $D=16
M72 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=42000 $Y=165550 $D=16
M73 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=44400 $Y=165550 $D=16
M74 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=97085 $D=16
M75 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=101995 $D=16
M76 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=103565 $D=16
M77 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=108475 $D=16
M78 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=110045 $D=16
M79 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=114955 $D=16
M80 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=116525 $D=16
M81 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=121435 $D=16
M82 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=123005 $D=16
M83 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=127915 $D=16
M84 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=59400 $Y=165550 $D=16
M85 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=61800 $Y=165550 $D=16
M86 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=64200 $Y=165550 $D=16
M87 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=66600 $Y=165550 $D=16
M88 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=69000 $Y=165550 $D=16
M89 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=71400 $Y=165550 $D=16
M90 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=73800 $Y=165550 $D=16
M91 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=76200 $Y=165550 $D=16
M92 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=78600 $Y=165550 $D=16
M93 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=81000 $Y=165550 $D=16
M94 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=83400 $Y=165550 $D=16
M95 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=85800 $Y=165550 $D=16
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4
** N=6 EP=4 IP=6 FDC=96
X0 1 4 2 3 pad_in $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_67
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_66
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_65
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_64
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_63
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pad_corner
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_32
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_16
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_8
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_2
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_01
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_62
** N=4 EP=0 IP=44 FDC=0
.ENDS
***************************************
.SUBCKT pad_fill_005
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_61
** N=4 EP=0 IP=72 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_59
** N=5 EP=0 IP=72 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57
** N=4 EP=0 IP=72 FDC=0
.ENDS
***************************************
.SUBCKT ICV_56
** N=4 EP=0 IP=40 FDC=0
.ENDS
***************************************
.SUBCKT ICV_55
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_60
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_58
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1 VSS VDD
** N=38 EP=2 IP=1 FDC=1
D0 VSS VDD pdio_m AREA=9e-10 PJ=0.00012 $X=8570 $Y=96300 $D=31
.ENDS
***************************************
.SUBCKT ICV_4 1 2 4
** N=7 EP=3 IP=6 FDC=96
X0 1 4 2 7 pad_in $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_54
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT bridge_soc_top_VIA15
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_53
** N=6 EP=0 IP=73 FDC=0
.ENDS
***************************************
.SUBCKT FILL2
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFFQSRX1 D CLK SETB RESETB VSS VDD Q
** N=34 EP=7 IP=0 FDC=40
M0 VSS D 20 VSS N L=1.8e-07 W=2.2e-07 $X=945 $Y=750 $D=0
M1 10 CLK VSS VSS N L=1.8e-07 W=2.2e-07 $X=1745 $Y=750 $D=0
M2 11 10 20 VSS N L=1.8e-07 W=2.2e-07 $X=3245 $Y=755 $D=0
M3 12 11 VSS VSS N L=1.8e-07 W=2.2e-07 $X=4745 $Y=755 $D=0
M4 13 12 VSS VSS N L=1.8e-07 W=2.2e-07 $X=6250 $Y=760 $D=0
M5 VSS 14 13 VSS N L=1.8e-07 W=2.2e-07 $X=7050 $Y=760 $D=0
M6 15 13 VSS VSS N L=1.8e-07 W=2.2e-07 $X=7850 $Y=1120 $D=0
M7 VSS SETB 14 VSS N L=1.8e-07 W=2.2e-07 $X=9355 $Y=755 $D=0
M8 22 CLK 11 VSS N L=1.8e-07 W=2.2e-07 $X=10860 $Y=750 $D=0
M9 33 15 VSS VSS N L=1.8e-07 W=4.4e-07 $X=12320 $Y=965 $D=0
M10 22 RESETB 33 VSS N L=1.8e-07 W=4.4e-07 $X=13040 $Y=965 $D=0
M11 16 CLK 15 VSS N L=1.8e-07 W=2.2e-07 $X=14500 $Y=755 $D=0
M12 34 16 VSS VSS N L=1.8e-07 W=4.4e-07 $X=15960 $Y=740 $D=0
M13 17 RESETB 34 VSS N L=1.8e-07 W=4.4e-07 $X=16680 $Y=740 $D=0
M14 18 17 VSS VSS N L=1.8e-07 W=2.2e-07 $X=18140 $Y=755 $D=0
M15 19 18 VSS VSS N L=1.8e-07 W=2.2e-07 $X=19640 $Y=755 $D=0
M16 VSS 14 19 VSS N L=1.8e-07 W=2.2e-07 $X=20440 $Y=755 $D=0
M17 24 19 VSS VSS N L=1.8e-07 W=2.2e-07 $X=21240 $Y=755 $D=0
M18 16 10 24 VSS N L=1.8e-07 W=2.2e-07 $X=22740 $Y=755 $D=0
M19 Q 17 VSS VSS N L=1.8e-07 W=2.2e-07 $X=24240 $Y=755 $D=0
M20 VDD D 20 VDD P L=1.8e-07 W=4.4e-07 $X=945 $Y=2705 $D=16
M21 10 CLK VDD VDD P L=1.8e-07 W=4.4e-07 $X=1665 $Y=2705 $D=16
M22 11 CLK 20 VDD P L=1.8e-07 W=4.4e-07 $X=3245 $Y=2725 $D=16
M23 12 11 VDD VDD P L=1.8e-07 W=4.4e-07 $X=4745 $Y=2725 $D=16
M24 21 12 13 VDD P L=1.8e-07 W=8.8e-07 $X=6250 $Y=2300 $D=16
M25 VDD 14 21 VDD P L=1.8e-07 W=8.8e-07 $X=6970 $Y=2300 $D=16
M26 15 13 VDD VDD P L=1.8e-07 W=4.4e-07 $X=7730 $Y=2520 $D=16
M27 VDD SETB 14 VDD P L=1.8e-07 W=4.4e-07 $X=9355 $Y=2535 $D=16
M28 22 10 11 VDD P L=1.8e-07 W=4.4e-07 $X=10815 $Y=2505 $D=16
M29 22 15 VDD VDD P L=1.8e-07 W=4.4e-07 $X=12320 $Y=2505 $D=16
M30 VDD RESETB 22 VDD P L=1.8e-07 W=4.4e-07 $X=13040 $Y=2505 $D=16
M31 16 10 15 VDD P L=1.8e-07 W=4.4e-07 $X=14500 $Y=2505 $D=16
M32 17 16 VDD VDD P L=1.8e-07 W=4.4e-07 $X=15960 $Y=2665 $D=16
M33 VDD RESETB 17 VDD P L=1.8e-07 W=4.4e-07 $X=16680 $Y=2665 $D=16
M34 18 17 VDD VDD P L=1.8e-07 W=4.4e-07 $X=18140 $Y=2725 $D=16
M35 23 18 19 VDD P L=1.8e-07 W=8.8e-07 $X=19640 $Y=2285 $D=16
M36 VDD 14 23 VDD P L=1.8e-07 W=8.8e-07 $X=20360 $Y=2285 $D=16
M37 24 19 VDD VDD P L=1.8e-07 W=4.4e-07 $X=21120 $Y=2505 $D=16
M38 16 CLK 24 VDD P L=1.8e-07 W=4.4e-07 $X=22740 $Y=2505 $D=16
M39 Q 17 VDD VDD P L=1.8e-07 W=4.4e-07 $X=24200 $Y=2505 $D=16
.ENDS
***************************************
.SUBCKT FILL32
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_43
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT FILL16
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL4
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2X1 A B VSS VDD Z
** N=9 EP=5 IP=0 FDC=4
M0 9 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=985 $Y=745 $D=0
M1 Z B 9 VSS N L=1.8e-07 W=4.4e-07 $X=1705 $Y=745 $D=0
M2 Z A VDD VDD P L=1.8e-07 W=4.4e-07 $X=985 $Y=2670 $D=16
M3 VDD B Z VDD P L=1.8e-07 W=4.4e-07 $X=1705 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT FILL8
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL1
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2X1 A B VSS VDD Z
** N=10 EP=5 IP=0 FDC=6
M0 10 A 8 VSS N L=1.8e-07 W=4.4e-07 $X=905 $Y=750 $D=0
M1 VSS B 10 VSS N L=1.8e-07 W=4.4e-07 $X=1625 $Y=750 $D=0
M2 Z 8 VSS VSS N L=1.8e-07 W=2.2e-07 $X=2385 $Y=860 $D=0
M3 8 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=905 $Y=2670 $D=16
M4 VDD B 8 VDD P L=1.8e-07 W=4.4e-07 $X=1625 $Y=2670 $D=16
M5 Z 8 VDD VDD P L=1.8e-07 W=4.4e-07 $X=2385 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT MUX2X1 A S B VSS VDD Z
** N=16 EP=6 IP=0 FDC=12
M0 VSS S 9 VSS N L=1.8e-07 W=4.4e-07 $X=940 $Y=960 $D=0
M1 15 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=1660 $Y=960 $D=0
M2 10 9 15 VSS N L=1.8e-07 W=4.4e-07 $X=2380 $Y=960 $D=0
M3 16 S 10 VSS N L=1.8e-07 W=4.4e-07 $X=3100 $Y=960 $D=0
M4 VSS B 16 VSS N L=1.8e-07 W=4.4e-07 $X=3920 $Y=740 $D=0
M5 Z 10 VSS VSS N L=1.8e-07 W=4.4e-07 $X=4640 $Y=740 $D=0
M6 VDD S 9 VDD P L=1.8e-07 W=4.4e-07 $X=940 $Y=2520 $D=16
M7 11 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1660 $Y=2520 $D=16
M8 10 S 11 VDD P L=1.8e-07 W=4.4e-07 $X=2380 $Y=2520 $D=16
M9 12 9 10 VDD P L=1.8e-07 W=4.4e-07 $X=3100 $Y=2520 $D=16
M10 VDD B 12 VDD P L=1.8e-07 W=4.4e-07 $X=3920 $Y=2735 $D=16
M11 Z 10 VDD VDD P L=1.8e-07 W=4.4e-07 $X=4640 $Y=2735 $D=16
.ENDS
***************************************
.SUBCKT NOR2X1 A B VSS VDD Z
** N=10 EP=5 IP=0 FDC=4
M0 Z A VSS VSS N L=1.8e-07 W=2.2e-07 $X=925 $Y=760 $D=0
M1 VSS B Z VSS N L=1.8e-07 W=2.2e-07 $X=1725 $Y=760 $D=0
M2 8 A VDD VDD P L=1.8e-07 W=8.8e-07 $X=925 $Y=2300 $D=16
M3 Z B 8 VDD P L=1.8e-07 W=8.8e-07 $X=1645 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT INVX2 A VSS VDD Z
** N=6 EP=4 IP=0 FDC=2
M0 Z A VSS VSS N L=1.8e-07 W=4.4e-07 $X=740 $Y=740 $D=0
M1 Z A VDD VDD P L=1.8e-07 W=8.8e-07 $X=740 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT ICV_52 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 29
** N=40 EP=28 IP=371 FDC=298
X13 25 24 2 23 1 2 3 DFFQSRX1 $T=339600 317200 0 180 $X=313970 $Y=312645
X14 26 24 2 23 1 2 4 DFFQSRX1 $T=339600 317200 1 180 $X=313970 $Y=316810
X15 27 24 2 23 1 2 5 DFFQSRX1 $T=339600 325040 0 180 $X=313970 $Y=320485
X16 33 24 23 2 1 2 16 DFFQSRX1 $T=619600 317200 1 0 $X=619170 $Y=312645
X17 37 24 23 2 1 2 18 DFFQSRX1 $T=619600 317200 0 0 $X=619170 $Y=316810
X18 29 24 23 2 1 2 21 DFFQSRX1 $T=619600 325040 1 0 $X=619170 $Y=320485
X60 6 3 1 2 7 NAND2X1 $T=387760 325040 1 0 $X=387330 $Y=320485
X61 8 9 1 2 32 NAND2X1 $T=425840 325040 1 0 $X=425410 $Y=320485
X62 32 11 1 2 10 NAND2X1 $T=431440 325040 1 0 $X=431010 $Y=320485
X69 14 13 1 2 12 AND2X1 $T=449920 325040 0 180 $X=446130 $Y=320485
X70 34 15 1 2 33 AND2X1 $T=583200 325040 0 180 $X=579410 $Y=320485
X71 18 16 1 2 19 AND2X1 $T=598320 317200 0 0 $X=597890 $Y=316810
X72 20 15 1 2 37 AND2X1 $T=603920 317200 0 0 $X=603490 $Y=316810
X73 35 17 16 1 2 34 MUX2X1 $T=591040 325040 0 180 $X=585010 $Y=320485
X74 16 18 1 2 36 NOR2X1 $T=594400 317200 1 180 $X=591170 $Y=316810
X75 36 19 1 2 35 NOR2X1 $T=595520 317200 0 0 $X=595090 $Y=316810
X76 22 1 2 23 INVX2 $T=644800 317200 1 0 $X=644370 $Y=312645
.ENDS
***************************************
.SUBCKT ICV_44
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_41
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_49
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_50 1 2 3 4 5
** N=7 EP=5 IP=11 FDC=4
X0 3 4 1 2 5 NAND2X1 $T=1680 0 0 0 $X=1250 $Y=-390
.ENDS
***************************************
.SUBCKT ICV_37
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT NAND3X1 A B C VSS VDD Z
** N=10 EP=6 IP=0 FDC=6
M0 9 A VSS VSS N L=1.8e-07 W=6.6e-07 $X=1210 $Y=745 $D=0
M1 10 B 9 VSS N L=1.8e-07 W=6.6e-07 $X=1930 $Y=745 $D=0
M2 Z C 10 VSS N L=1.8e-07 W=6.6e-07 $X=2650 $Y=745 $D=0
M3 Z A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1210 $Y=2670 $D=16
M4 VDD B Z VDD P L=1.8e-07 W=4.4e-07 $X=1930 $Y=2670 $D=16
M5 Z C VDD VDD P L=1.8e-07 W=4.4e-07 $X=2650 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT ICV_42
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_48
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT OR2X1 A B VSS VDD Z
** N=12 EP=5 IP=0 FDC=6
M0 8 A VSS VSS N L=1.8e-07 W=2.2e-07 $X=835 $Y=760 $D=0
M1 VSS B 8 VSS N L=1.8e-07 W=2.2e-07 $X=1635 $Y=760 $D=0
M2 Z 8 VSS VSS N L=1.8e-07 W=2.2e-07 $X=2435 $Y=760 $D=0
M3 9 A 8 VDD P L=1.8e-07 W=8.8e-07 $X=835 $Y=2300 $D=16
M4 VDD B 9 VDD P L=1.8e-07 W=8.8e-07 $X=1555 $Y=2300 $D=16
M5 Z 8 VDD VDD P L=1.8e-07 W=4.4e-07 $X=2315 $Y=2520 $D=16
.ENDS
***************************************
.SUBCKT INVX8 A VSS VDD Z
** N=6 EP=4 IP=0 FDC=8
M0 Z A VSS VSS N L=1.8e-07 W=4.4e-07 $X=740 $Y=760 $D=0
M1 VSS A Z VSS N L=1.8e-07 W=4.4e-07 $X=1460 $Y=760 $D=0
M2 Z A VSS VSS N L=1.8e-07 W=4.4e-07 $X=2180 $Y=760 $D=0
M3 VSS A Z VSS N L=1.8e-07 W=4.4e-07 $X=2900 $Y=760 $D=0
M4 Z A VDD VDD P L=1.8e-07 W=8.8e-07 $X=740 $Y=2300 $D=16
M5 VDD A Z VDD P L=1.8e-07 W=8.8e-07 $X=1460 $Y=2300 $D=16
M6 Z A VDD VDD P L=1.8e-07 W=8.8e-07 $X=2180 $Y=2300 $D=16
M7 VDD A Z VDD P L=1.8e-07 W=8.8e-07 $X=2900 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT ANTENNA VSS A
** N=5 EP=2 IP=0 FDC=1
*.CALIBRE ISOLATED NETS: VDD
D0 VSS A DN AREA=3.9e-13 PJ=2.54e-06 $X=300 $Y=655 $D=26
.ENDS
***************************************
.SUBCKT XOR2X1 B A VDD VSS Z
** N=11 EP=5 IP=0 FDC=10
M0 VSS B 10 VSS N L=1.8e-07 W=4.4e-07 $X=630 $Y=985 $D=0
M1 8 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=1350 $Y=985 $D=0
M2 9 8 10 VSS N L=1.8e-07 W=4.4e-07 $X=3205 $Y=1000 $D=0
M3 B A 9 VSS N L=1.8e-07 W=4.4e-07 $X=3925 $Y=1000 $D=0
M4 Z 9 VSS VSS N L=1.8e-07 W=4.4e-07 $X=5345 $Y=1000 $D=0
M5 VDD B 10 VDD P L=1.8e-07 W=4.4e-07 $X=630 $Y=2435 $D=16
M6 8 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1350 $Y=2435 $D=16
M7 9 A 10 VDD P L=1.8e-07 W=4.4e-07 $X=3205 $Y=2435 $D=16
M8 B 8 9 VDD P L=1.8e-07 W=4.4e-07 $X=3925 $Y=2435 $D=16
M9 Z 9 VDD VDD P L=1.8e-07 W=4.4e-07 $X=5345 $Y=2435 $D=16
.ENDS
***************************************
.SUBCKT ICV_51 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94
** N=510 EP=94 IP=5567 FDC=6194
M0 97 1 2 2 N L=1.8e-07 W=4.4e-07 $X=419790 $Y=396360 $D=0
M1 2 1 97 2 N L=1.8e-07 W=4.4e-07 $X=420510 $Y=396360 $D=0
M2 97 1 3 3 P L=1.8e-07 W=8.8e-07 $X=419790 $Y=397900 $D=16
M3 3 1 97 3 P L=1.8e-07 W=8.8e-07 $X=420510 $Y=397900 $D=16
X47 193 82 3 83 2 3 102 DFFQSRX1 $T=314400 325040 0 0 $X=313970 $Y=324650
X48 131 82 83 3 2 3 103 DFFQSRX1 $T=314400 332880 1 0 $X=313970 $Y=328325
X49 170 82 3 83 2 3 98 DFFQSRX1 $T=339600 340720 0 180 $X=313970 $Y=336165
X50 188 82 3 83 2 3 104 DFFQSRX1 $T=314400 340720 0 0 $X=313970 $Y=340330
X51 183 82 3 83 2 3 105 DFFQSRX1 $T=314400 356400 0 0 $X=313970 $Y=356010
X52 126 82 83 3 2 3 106 DFFQSRX1 $T=314400 364240 1 0 $X=313970 $Y=359685
X53 134 82 83 3 2 3 107 DFFQSRX1 $T=314400 411280 0 0 $X=313970 $Y=410890
X54 3 82 3 83 2 3 4 DFFQSRX1 $T=349120 403440 1 180 $X=323490 $Y=403050
X55 101 82 83 3 2 3 5 DFFQSRX1 $T=353600 411280 0 180 $X=327970 $Y=406725
X56 129 82 83 3 2 3 99 DFFQSRX1 $T=355280 387760 0 180 $X=329650 $Y=383205
X57 110 82 83 3 2 3 100 DFFQSRX1 $T=355840 379920 1 180 $X=330210 $Y=379530
X58 120 82 83 3 2 3 125 DFFQSRX1 $T=341840 348560 1 0 $X=341410 $Y=344005
X59 113 82 83 3 2 3 111 DFFQSRX1 $T=341840 348560 0 0 $X=341410 $Y=348170
X60 117 82 83 3 2 3 121 DFFQSRX1 $T=341840 372080 0 0 $X=341410 $Y=371690
X61 155 82 83 3 2 3 152 DFFQSRX1 $T=345200 372080 1 0 $X=344770 $Y=367525
X62 84 82 83 3 2 3 9 DFFQSRX1 $T=370400 426960 1 180 $X=344770 $Y=426570
X63 141 82 83 3 2 3 127 DFFQSRX1 $T=349120 403440 0 0 $X=348690 $Y=403050
X64 147 82 83 3 2 3 136 DFFQSRX1 $T=381040 379920 1 180 $X=355410 $Y=379530
X65 164 82 83 3 2 3 143 DFFQSRX1 $T=386640 387760 0 180 $X=361010 $Y=383205
X66 167 82 83 3 2 3 11 DFFQSRX1 $T=386640 411280 0 180 $X=361010 $Y=406725
X67 177 82 3 83 2 3 159 DFFQSRX1 $T=397280 348560 0 180 $X=371650 $Y=344005
X68 144 82 83 3 2 3 150 DFFQSRX1 $T=372080 348560 0 0 $X=371650 $Y=348170
X69 151 82 3 83 2 3 168 DFFQSRX1 $T=372080 372080 1 0 $X=371650 $Y=367525
X70 165 82 3 83 2 3 160 DFFQSRX1 $T=397280 372080 1 180 $X=371650 $Y=371690
X71 85 82 83 3 2 3 20 DFFQSRX1 $T=372080 426960 1 0 $X=371650 $Y=422405
X72 86 82 83 3 2 3 21 DFFQSRX1 $T=372080 426960 0 0 $X=371650 $Y=426570
X73 175 82 83 3 2 3 179 DFFQSRX1 $T=381040 379920 0 0 $X=380610 $Y=379530
X74 184 82 83 3 2 3 194 DFFQSRX1 $T=381600 403440 0 0 $X=381170 $Y=403050
X75 197 82 83 3 2 3 181 DFFQSRX1 $T=416880 387760 0 180 $X=391250 $Y=383205
X76 192 82 83 3 2 3 182 DFFQSRX1 $T=416880 411280 0 180 $X=391250 $Y=406725
X77 88 82 83 3 2 3 25 DFFQSRX1 $T=402320 426960 1 0 $X=401890 $Y=422405
X78 87 82 83 3 2 3 29 DFFQSRX1 $T=402320 426960 0 0 $X=401890 $Y=426570
X79 224 82 83 3 2 3 206 DFFQSRX1 $T=404000 372080 1 0 $X=403570 $Y=367525
X80 217 82 83 3 2 3 221 DFFQSRX1 $T=405680 348560 1 0 $X=405250 $Y=344005
X81 89 82 83 3 2 3 27 DFFQSRX1 $T=405680 348560 0 0 $X=405250 $Y=348170
X82 218 82 83 3 2 3 162 DFFQSRX1 $T=430880 372080 1 180 $X=405250 $Y=371690
X83 203 82 83 3 2 3 202 DFFQSRX1 $T=406240 379920 0 0 $X=405810 $Y=379530
X84 220 82 83 3 2 3 228 DFFQSRX1 $T=409040 403440 0 0 $X=408610 $Y=403050
X85 219 82 83 3 2 3 212 DFFQSRX1 $T=442080 411280 0 180 $X=416450 $Y=406725
X86 262 82 83 3 2 3 239 DFFQSRX1 $T=458320 348560 1 180 $X=432690 $Y=348170
X87 259 82 83 3 2 3 248 DFFQSRX1 $T=458320 372080 0 180 $X=432690 $Y=367525
X88 243 82 83 3 2 3 254 DFFQSRX1 $T=433120 372080 0 0 $X=432690 $Y=371690
X89 270 82 83 3 2 3 32 DFFQSRX1 $T=458320 426960 0 180 $X=432690 $Y=422405
X90 90 82 83 3 2 3 33 DFFQSRX1 $T=458320 426960 1 180 $X=432690 $Y=426570
X91 267 82 83 3 2 3 253 DFFQSRX1 $T=461680 348560 0 180 $X=436050 $Y=344005
X92 263 82 83 3 2 3 272 DFFQSRX1 $T=437040 379920 0 0 $X=436610 $Y=379530
X93 269 82 83 3 2 3 251 DFFQSRX1 $T=438160 387760 1 0 $X=437730 $Y=383205
X94 261 82 83 3 2 3 266 DFFQSRX1 $T=442080 411280 1 0 $X=441650 $Y=406725
X95 275 82 83 3 2 3 271 DFFQSRX1 $T=477360 403440 1 180 $X=451730 $Y=403050
X96 260 82 83 3 2 3 36 DFFQSRX1 $T=488560 348560 1 180 $X=462930 $Y=348170
X97 277 82 83 3 2 3 287 DFFQSRX1 $T=463360 372080 0 0 $X=462930 $Y=371690
X98 281 82 83 3 2 3 288 DFFQSRX1 $T=463360 426960 0 0 $X=462930 $Y=426570
X99 295 82 83 3 2 3 314 DFFQSRX1 $T=466720 348560 1 0 $X=466290 $Y=344005
X100 306 82 83 3 2 3 283 DFFQSRX1 $T=491920 372080 0 180 $X=466290 $Y=367525
X101 91 82 83 3 2 3 282 DFFQSRX1 $T=491920 426960 0 180 $X=466290 $Y=422405
X102 308 82 83 3 2 3 298 DFFQSRX1 $T=506480 387760 0 180 $X=480850 $Y=383205
X103 315 82 83 3 2 3 297 DFFQSRX1 $T=506480 403440 1 180 $X=480850 $Y=403050
X104 322 82 83 3 2 3 303 DFFQSRX1 $T=508160 379920 1 180 $X=482530 $Y=379530
X105 326 82 83 3 2 3 304 DFFQSRX1 $T=508160 411280 0 180 $X=482530 $Y=406725
X106 311 82 83 3 2 3 324 DFFQSRX1 $T=493600 348560 1 0 $X=493170 $Y=344005
X107 317 82 83 3 2 3 327 DFFQSRX1 $T=493600 348560 0 0 $X=493170 $Y=348170
X108 331 82 83 3 2 3 330 DFFQSRX1 $T=493600 372080 1 0 $X=493170 $Y=367525
X109 323 82 83 3 2 3 54 DFFQSRX1 $T=493600 426960 1 0 $X=493170 $Y=422405
X110 301 82 83 3 2 3 292 DFFQSRX1 $T=493600 426960 0 0 $X=493170 $Y=426570
X111 372 82 83 3 2 3 320 DFFQSRX1 $T=522160 372080 1 180 $X=496530 $Y=371690
X112 354 82 83 3 2 3 338 DFFQSRX1 $T=538400 379920 1 180 $X=512770 $Y=379530
X113 364 82 83 3 2 3 339 DFFQSRX1 $T=538400 387760 0 180 $X=512770 $Y=383205
X114 366 82 83 3 2 3 340 DFFQSRX1 $T=538400 403440 1 180 $X=512770 $Y=403050
X115 347 82 83 3 2 3 341 DFFQSRX1 $T=538400 411280 0 180 $X=512770 $Y=406725
X116 334 82 83 3 2 3 346 DFFQSRX1 $T=524400 348560 1 0 $X=523970 $Y=344005
X117 337 82 83 3 2 3 343 DFFQSRX1 $T=524400 348560 0 0 $X=523970 $Y=348170
X118 370 82 83 3 2 3 352 DFFQSRX1 $T=549600 372080 0 180 $X=523970 $Y=367525
X119 373 82 83 3 2 3 360 DFFQSRX1 $T=549600 372080 1 180 $X=523970 $Y=371690
X120 92 82 83 3 2 3 57 DFFQSRX1 $T=549600 426960 0 180 $X=523970 $Y=422405
X121 285 82 83 3 2 3 49 DFFQSRX1 $T=524400 426960 0 0 $X=523970 $Y=426570
X122 374 82 83 3 2 3 357 DFFQSRX1 $T=563600 379920 1 180 $X=537970 $Y=379530
X123 290 82 83 3 2 3 305 DFFQSRX1 $T=563600 387760 0 180 $X=537970 $Y=383205
X124 369 82 83 3 2 3 61 DFFQSRX1 $T=563600 403440 1 180 $X=537970 $Y=403050
X125 382 82 83 3 2 3 387 DFFQSRX1 $T=558000 348560 1 0 $X=557570 $Y=344005
X126 419 82 3 83 2 3 388 DFFQSRX1 $T=558000 348560 0 0 $X=557570 $Y=348170
X127 389 82 3 83 2 3 390 DFFQSRX1 $T=558000 372080 1 0 $X=557570 $Y=367525
X128 413 82 3 83 2 3 391 DFFQSRX1 $T=558000 372080 0 0 $X=557570 $Y=371690
X129 399 82 83 3 2 3 375 DFFQSRX1 $T=583200 426960 0 180 $X=557570 $Y=422405
X130 62 82 83 3 2 3 376 DFFQSRX1 $T=592160 379920 1 180 $X=566530 $Y=379530
X131 398 82 83 3 2 3 377 DFFQSRX1 $T=593840 411280 0 180 $X=568210 $Y=406725
X132 397 82 83 3 2 3 378 DFFQSRX1 $T=594400 403440 1 180 $X=568770 $Y=403050
X133 417 82 83 3 2 3 379 DFFQSRX1 $T=599440 387760 0 180 $X=573810 $Y=383205
X134 386 82 83 3 2 3 403 DFFQSRX1 $T=584880 348560 1 0 $X=584450 $Y=344005
X135 393 82 3 83 2 3 410 DFFQSRX1 $T=584880 348560 0 0 $X=584450 $Y=348170
X136 93 82 83 3 2 3 71 DFFQSRX1 $T=584880 426960 1 0 $X=584450 $Y=422405
X137 94 82 83 3 2 3 67 DFFQSRX1 $T=613440 426960 1 180 $X=587810 $Y=426570
X138 435 82 3 83 2 3 426 DFFQSRX1 $T=592720 379920 0 0 $X=592290 $Y=379530
X139 428 82 83 3 2 3 432 DFFQSRX1 $T=594400 403440 0 0 $X=593970 $Y=403050
X140 461 82 83 3 2 3 429 DFFQSRX1 $T=627440 411280 0 180 $X=601810 $Y=406725
X141 471 82 83 3 2 3 434 DFFQSRX1 $T=629680 387760 0 180 $X=604050 $Y=383205
X142 474 82 3 83 2 3 454 DFFQSRX1 $T=640880 348560 0 180 $X=615250 $Y=344005
X143 460 82 3 83 2 3 450 DFFQSRX1 $T=640880 372080 1 180 $X=615250 $Y=371690
X144 475 82 83 3 2 3 76 DFFQSRX1 $T=640880 426960 1 180 $X=615250 $Y=426570
X145 439 82 83 3 2 3 412 DFFQSRX1 $T=619600 332880 1 0 $X=619170 $Y=328325
X146 456 82 3 83 2 3 451 DFFQSRX1 $T=619600 340720 1 0 $X=619170 $Y=336165
X147 470 82 3 83 2 3 444 DFFQSRX1 $T=619600 356400 1 0 $X=619170 $Y=351845
X148 463 82 3 83 2 3 442 DFFQSRX1 $T=619600 364240 0 0 $X=619170 $Y=363850
X149 462 82 83 3 2 3 455 DFFQSRX1 $T=619600 395600 1 0 $X=619170 $Y=391045
X150 468 82 83 3 2 3 464 DFFQSRX1 $T=619600 403440 0 0 $X=619170 $Y=403050
X151 478 82 83 3 2 3 481 DFFQSRX1 $T=625200 403440 1 0 $X=624770 $Y=398885
X152 482 82 83 3 2 3 472 DFFQSRX1 $T=650960 372080 0 180 $X=625330 $Y=367525
X153 484 82 83 3 2 3 473 DFFQSRX1 $T=652080 426960 0 180 $X=626450 $Y=422405
X154 479 82 83 3 2 3 480 DFFQSRX1 $T=627440 419120 1 0 $X=627010 $Y=414565
X155 3 82 3 83 2 3 81 DFFQSRX1 $T=629120 325040 0 0 $X=628690 $Y=324650
X156 483 82 83 3 2 3 477 DFFQSRX1 $T=654880 387760 0 180 $X=629250 $Y=383205
X326 7 111 2 3 109 NAND2X1 $T=339040 348560 0 0 $X=338610 $Y=348170
X327 108 112 2 3 110 NAND2X1 $T=339040 372080 1 0 $X=338610 $Y=367525
X328 109 115 2 3 113 NAND2X1 $T=341280 356400 1 0 $X=340850 $Y=351845
X329 7 100 2 3 108 NAND2X1 $T=341840 372080 1 0 $X=341410 $Y=367525
X330 7 121 2 3 114 NAND2X1 $T=342400 379920 1 0 $X=341970 $Y=375365
X331 118 123 2 3 120 NAND2X1 $T=342960 340720 0 0 $X=342530 $Y=340330
X332 7 99 2 3 122 NAND2X1 $T=342960 395600 0 0 $X=342530 $Y=395210
X333 10 106 2 3 115 NAND2X1 $T=347440 356400 0 180 $X=344210 $Y=351845
X334 10 100 2 3 124 NAND2X1 $T=345200 364240 0 0 $X=344770 $Y=363850
X335 7 125 2 3 118 NAND2X1 $T=346320 340720 0 0 $X=345890 $Y=340330
X336 10 111 2 3 123 NAND2X1 $T=350240 356400 0 180 $X=347010 $Y=351845
X337 116 124 2 3 126 NAND2X1 $T=348000 364240 0 0 $X=347570 $Y=363850
X338 10 99 2 3 119 NAND2X1 $T=351360 387760 1 180 $X=348130 $Y=387370
X339 122 128 2 3 129 NAND2X1 $T=349120 395600 0 0 $X=348690 $Y=395210
X340 10 127 2 3 128 NAND2X1 $T=351920 403440 0 180 $X=348690 $Y=398885
X341 10 121 2 3 112 NAND2X1 $T=350800 364240 0 0 $X=350370 $Y=363850
X342 132 130 2 3 131 NAND2X1 $T=354160 340720 1 180 $X=350930 $Y=340330
X343 7 107 2 3 133 NAND2X1 $T=355840 411280 1 180 $X=352610 $Y=410890
X344 7 127 2 3 137 NAND2X1 $T=354720 403440 1 0 $X=354290 $Y=398885
X345 10 103 2 3 138 NAND2X1 $T=355280 356400 1 0 $X=354850 $Y=351845
X346 10 107 2 3 140 NAND2X1 $T=361440 411280 1 180 $X=358210 $Y=410890
X347 10 9 2 3 139 NAND2X1 $T=359200 419120 0 0 $X=358770 $Y=418730
X348 145 138 2 3 144 NAND2X1 $T=364240 356400 0 180 $X=361010 $Y=351845
X349 7 150 2 3 145 NAND2X1 $T=367040 356400 1 0 $X=366610 $Y=351845
X350 10 150 2 3 148 NAND2X1 $T=367040 364240 1 0 $X=366610 $Y=359685
X351 158 148 2 3 155 NAND2X1 $T=372640 364240 0 180 $X=369410 $Y=359685
X352 160 162 2 3 156 NAND2X1 $T=372080 332880 1 0 $X=371650 $Y=328325
X353 7 152 2 3 158 NAND2X1 $T=373200 364240 1 0 $X=372770 $Y=359685
X354 16 14 2 3 163 NAND2X1 $T=382720 325040 1 180 $X=379490 $Y=324650
X355 10 152 2 3 171 NAND2X1 $T=383840 364240 0 180 $X=380610 $Y=359685
X356 168 162 2 3 172 NAND2X1 $T=381600 356400 1 0 $X=381170 $Y=351845
X357 16 159 2 3 173 NAND2X1 $T=387760 332880 0 180 $X=384530 $Y=328325
X358 1 5 2 3 142 NAND2X1 $T=389440 419120 1 180 $X=386210 $Y=418730
X359 97 13 2 3 153 NAND2X1 $T=390000 356400 0 180 $X=386770 $Y=351845
X360 1 15 2 3 135 NAND2X1 $T=392240 419120 1 180 $X=389010 $Y=418730
X361 16 105 2 3 180 NAND2X1 $T=390000 356400 1 0 $X=389570 $Y=351845
X362 7 21 2 3 23 NAND2X1 $T=400080 426960 1 180 $X=396850 $Y=426570
X363 22 162 2 3 186 NAND2X1 $T=397840 325040 0 0 $X=397410 $Y=324650
X364 104 162 2 3 189 NAND2X1 $T=400640 340720 0 180 $X=397410 $Y=336165
X365 194 162 2 3 187 NAND2X1 $T=402320 356400 0 180 $X=399090 $Y=351845
X366 190 194 2 3 185 NAND2X1 $T=399520 364240 1 0 $X=399090 $Y=359685
X367 16 22 2 3 195 NAND2X1 $T=403440 325040 1 180 $X=400210 $Y=324650
X368 16 104 2 3 191 NAND2X1 $T=405680 348560 1 180 $X=402450 $Y=348170
X369 102 162 2 3 198 NAND2X1 $T=407360 332880 0 180 $X=404130 $Y=328325
X370 181 202 2 3 205 NAND2X1 $T=414640 387760 1 180 $X=411410 $Y=387370
X371 162 206 2 3 13 NAND2X1 $T=415760 340720 1 180 $X=412530 $Y=340330
X372 209 210 2 3 211 NAND2X1 $T=414080 340720 1 0 $X=413650 $Y=336165
X373 211 162 2 3 213 NAND2X1 $T=416320 332880 1 0 $X=415890 $Y=328325
X374 190 205 2 3 207 NAND2X1 $T=419680 387760 0 180 $X=416450 $Y=383205
X375 223 208 2 3 218 NAND2X1 $T=420800 379920 0 180 $X=417570 $Y=375365
X376 222 210 2 3 226 NAND2X1 $T=420800 387760 1 0 $X=420370 $Y=383205
X377 226 190 2 3 229 NAND2X1 $T=423600 387760 1 0 $X=423170 $Y=383205
X378 231 210 2 3 230 NAND2X1 $T=427520 332880 1 180 $X=424290 $Y=332490
X379 214 221 2 3 231 NAND2X1 $T=424720 340720 0 0 $X=424290 $Y=340330
X380 1 182 2 3 28 NAND2X1 $T=427520 419120 1 180 $X=424290 $Y=418730
X381 230 162 2 3 232 NAND2X1 $T=425280 325040 0 0 $X=424850 $Y=324650
X382 235 162 2 3 234 NAND2X1 $T=429200 356400 1 180 $X=425970 $Y=356010
X383 238 162 2 3 236 NAND2X1 $T=429760 340720 0 180 $X=426530 $Y=336165
X384 210 240 2 3 235 NAND2X1 $T=427520 356400 1 0 $X=427090 $Y=351845
X385 97 245 2 3 243 NAND2X1 $T=430320 372080 1 0 $X=429890 $Y=367525
X386 1 228 2 3 31 NAND2X1 $T=433120 426960 0 180 $X=429890 $Y=422405
X387 241 249 2 3 233 NAND2X1 $T=431440 340720 0 0 $X=431010 $Y=340330
X388 234 239 2 3 247 NAND2X1 $T=431440 356400 0 0 $X=431010 $Y=356010
X389 26 244 2 3 34 NAND2X1 $T=435920 325040 1 180 $X=432690 $Y=324650
X390 1 212 2 3 35 NAND2X1 $T=433120 419120 1 0 $X=432690 $Y=414565
X391 7 32 2 3 252 NAND2X1 $T=434800 419120 0 0 $X=434370 $Y=418730
X392 10 246 2 3 257 NAND2X1 $T=440960 356400 1 180 $X=437730 $Y=356010
X393 257 247 2 3 262 NAND2X1 $T=446560 356400 1 180 $X=443330 $Y=356010
X394 10 254 2 3 264 NAND2X1 $T=447680 364240 0 0 $X=447250 $Y=363850
X395 190 272 2 3 265 NAND2X1 $T=450480 364240 0 0 $X=450050 $Y=363850
X396 10 272 2 3 273 NAND2X1 $T=453840 364240 0 0 $X=453410 $Y=363850
X397 1 266 2 3 268 NAND2X1 $T=461120 419120 0 180 $X=457890 $Y=414565
X398 1 39 2 3 41 NAND2X1 $T=461120 419120 1 180 $X=457890 $Y=418730
X399 1 43 2 3 42 NAND2X1 $T=458320 426960 1 0 $X=457890 $Y=422405
X400 190 271 2 3 274 NAND2X1 $T=458880 372080 1 0 $X=458450 $Y=367525
X401 10 271 2 3 276 NAND2X1 $T=461680 379920 1 0 $X=461250 $Y=375365
X402 190 288 2 3 286 NAND2X1 $T=469520 379920 1 0 $X=469090 $Y=375365
X403 190 50 2 3 284 NAND2X1 $T=470080 356400 0 0 $X=469650 $Y=356010
X404 289 291 2 3 290 NAND2X1 $T=474560 340720 1 0 $X=474130 $Y=336165
X405 10 288 2 3 278 NAND2X1 $T=475120 379920 1 0 $X=474690 $Y=375365
X406 10 50 2 3 291 NAND2X1 $T=479040 340720 1 180 $X=475810 $Y=340330
X407 10 292 2 3 279 NAND2X1 $T=479600 356400 1 180 $X=476370 $Y=356010
X408 10 287 2 3 293 NAND2X1 $T=477920 364240 1 0 $X=477490 $Y=359685
X409 7 297 2 3 299 NAND2X1 $T=482960 419120 0 180 $X=479730 $Y=414565
X410 302 300 2 3 301 NAND2X1 $T=484080 356400 0 180 $X=480850 $Y=351845
X411 10 283 2 3 300 NAND2X1 $T=481840 356400 0 0 $X=481410 $Y=356010
X412 10 305 2 3 296 NAND2X1 $T=482400 340720 0 0 $X=481970 $Y=340330
X413 10 297 2 3 51 NAND2X1 $T=485760 419120 0 180 $X=482530 $Y=414565
X414 7 282 2 3 52 NAND2X1 $T=483520 419120 0 0 $X=483090 $Y=418730
X415 7 305 2 3 289 NAND2X1 $T=486880 340720 0 180 $X=483650 $Y=336165
X416 307 293 2 3 306 NAND2X1 $T=488000 364240 0 180 $X=484770 $Y=359685
X417 7 283 2 3 307 NAND2X1 $T=488560 356400 1 180 $X=485330 $Y=356010
X418 7 292 2 3 302 NAND2X1 $T=489120 356400 0 180 $X=485890 $Y=351845
X419 1 48 2 3 309 NAND2X1 $T=489680 419120 0 180 $X=486450 $Y=414565
X420 10 282 2 3 312 NAND2X1 $T=492480 419120 0 180 $X=489250 $Y=414565
X421 1 49 2 3 53 NAND2X1 $T=493040 426960 1 180 $X=489810 $Y=426570
X422 10 314 2 3 313 NAND2X1 $T=497520 332880 1 180 $X=494290 $Y=332490
X423 319 316 2 3 317 NAND2X1 $T=497520 340720 1 180 $X=494290 $Y=340330
X424 1 298 2 3 318 NAND2X1 $T=494720 419120 1 0 $X=494290 $Y=414565
X425 1 303 2 3 321 NAND2X1 $T=495840 411280 0 0 $X=495410 $Y=410890
X426 10 324 2 3 316 NAND2X1 $T=497520 340720 0 0 $X=497090 $Y=340330
X427 7 324 2 3 310 NAND2X1 $T=502000 332880 1 180 $X=498770 $Y=332490
X428 7 327 2 3 319 NAND2X1 $T=500320 340720 0 0 $X=499890 $Y=340330
X429 7 304 2 3 328 NAND2X1 $T=502000 411280 0 0 $X=501570 $Y=410890
X430 329 332 2 3 331 NAND2X1 $T=504240 340720 0 0 $X=503810 $Y=340330
X431 10 330 2 3 333 NAND2X1 $T=510400 340720 0 180 $X=507170 $Y=336165
X432 10 304 2 3 55 NAND2X1 $T=507600 419120 1 0 $X=507170 $Y=414565
X433 335 333 2 3 334 NAND2X1 $T=511520 332880 1 180 $X=508290 $Y=332490
X434 10 327 2 3 332 NAND2X1 $T=509280 340720 0 0 $X=508850 $Y=340330
X435 1 57 2 3 56 NAND2X1 $T=509280 419120 0 0 $X=508850 $Y=418730
X436 336 342 2 3 337 NAND2X1 $T=511520 332880 0 0 $X=511090 $Y=332490
X437 7 343 2 3 336 NAND2X1 $T=513200 340720 1 0 $X=512770 $Y=336165
X438 10 58 2 3 325 NAND2X1 $T=513200 419120 0 0 $X=512770 $Y=418730
X439 10 339 2 3 345 NAND2X1 $T=518800 395600 0 180 $X=515570 $Y=391045
X440 10 346 2 3 342 NAND2X1 $T=519360 332880 1 180 $X=516130 $Y=332490
X441 7 346 2 3 335 NAND2X1 $T=519920 332880 0 180 $X=516690 $Y=328325
X442 10 320 2 3 348 NAND2X1 $T=518240 340720 1 0 $X=517810 $Y=336165
X443 10 59 2 3 344 NAND2X1 $T=518800 419120 0 0 $X=518370 $Y=418730
X444 7 339 2 3 351 NAND2X1 $T=522160 379920 0 180 $X=518930 $Y=375365
X445 10 352 2 3 353 NAND2X1 $T=523280 364240 0 180 $X=520050 $Y=359685
X446 355 353 2 3 354 NAND2X1 $T=523280 372080 0 180 $X=520050 $Y=367525
X447 7 340 2 3 356 NAND2X1 $T=523840 387760 1 180 $X=520610 $Y=387370
X448 10 357 2 3 359 NAND2X1 $T=524960 356400 1 180 $X=521730 $Y=356010
X449 10 338 2 3 358 NAND2X1 $T=522160 379920 1 0 $X=521730 $Y=375365
X450 10 343 2 3 361 NAND2X1 $T=523280 340720 1 0 $X=522850 $Y=336165
X451 10 360 2 3 362 NAND2X1 $T=526080 364240 0 180 $X=522850 $Y=359685
X452 7 341 2 3 349 NAND2X1 $T=523840 411280 0 0 $X=523410 $Y=410890
X453 7 61 2 3 363 NAND2X1 $T=524960 403440 1 0 $X=524530 $Y=398885
X454 351 358 2 3 364 NAND2X1 $T=528320 379920 0 180 $X=525090 $Y=375365
X455 7 320 2 3 365 NAND2X1 $T=528880 340720 0 180 $X=525650 $Y=336165
X456 356 345 2 3 366 NAND2X1 $T=528880 395600 0 180 $X=525650 $Y=391045
X457 7 357 2 3 367 NAND2X1 $T=530000 340720 1 180 $X=526770 $Y=340330
X458 7 360 2 3 368 NAND2X1 $T=530560 356400 1 180 $X=527330 $Y=356010
X459 371 362 2 3 370 NAND2X1 $T=530560 364240 0 180 $X=527330 $Y=359685
X460 363 350 2 3 369 NAND2X1 $T=530560 403440 0 180 $X=527330 $Y=398885
X461 7 338 2 3 355 NAND2X1 $T=528320 379920 1 0 $X=527890 $Y=375365
X462 365 361 2 3 372 NAND2X1 $T=531680 340720 0 180 $X=528450 $Y=336165
X463 368 359 2 3 373 NAND2X1 $T=533360 356400 1 180 $X=530130 $Y=356010
X464 7 352 2 3 371 NAND2X1 $T=533360 364240 0 180 $X=530130 $Y=359685
X465 367 348 2 3 374 NAND2X1 $T=534480 340720 0 180 $X=531250 $Y=336165
X466 381 377 2 3 380 NAND2X1 $T=580960 387760 1 180 $X=577730 $Y=387370
X467 381 376 2 3 384 NAND2X1 $T=583200 356400 0 180 $X=579970 $Y=351845
X468 381 378 2 3 383 NAND2X1 $T=583760 387760 1 180 $X=580530 $Y=387370
X469 403 390 2 3 404 NAND2X1 $T=587680 356400 0 0 $X=587250 $Y=356010
X470 403 410 2 3 407 NAND2X1 $T=594400 356400 0 180 $X=591170 $Y=351845
X471 412 391 2 3 401 NAND2X1 $T=594400 372080 0 180 $X=591170 $Y=367525
X472 381 379 2 3 409 NAND2X1 $T=594960 387760 1 180 $X=591730 $Y=387370
X473 412 390 2 3 411 NAND2X1 $T=596080 364240 0 180 $X=592850 $Y=359685
X474 403 391 2 3 416 NAND2X1 $T=597760 364240 1 180 $X=594530 $Y=363850
X475 381 432 2 3 431 NAND2X1 $T=601680 387760 1 0 $X=601250 $Y=383205
X476 63 420 2 3 425 NAND2X1 $T=606160 340720 1 180 $X=602930 $Y=340330
X477 403 426 2 3 433 NAND2X1 $T=606160 364240 1 180 $X=602930 $Y=363850
X478 68 421 2 3 439 NAND2X1 $T=608400 340720 0 180 $X=605170 $Y=336165
X479 403 442 2 3 438 NAND2X1 $T=605600 364240 1 0 $X=605170 $Y=359685
X480 412 403 2 3 63 NAND2X1 $T=610640 340720 1 180 $X=607410 $Y=340330
X481 412 444 2 3 436 NAND2X1 $T=607840 356400 0 0 $X=607410 $Y=356010
X482 412 450 2 3 440 NAND2X1 $T=609520 372080 0 0 $X=609090 $Y=371690
X483 412 454 2 3 449 NAND2X1 $T=610080 356400 1 0 $X=609650 $Y=351845
X484 381 455 2 3 458 NAND2X1 $T=616240 379920 0 180 $X=613010 $Y=375365
X485 403 454 2 3 459 NAND2X1 $T=614000 356400 1 0 $X=613570 $Y=351845
X486 403 444 2 3 452 NAND2X1 $T=614000 356400 0 0 $X=613570 $Y=356010
X487 403 450 2 3 453 NAND2X1 $T=620720 372080 0 180 $X=617490 $Y=367525
X488 381 434 2 3 466 NAND2X1 $T=619040 379920 0 0 $X=618610 $Y=379530
X489 412 451 2 3 465 NAND2X1 $T=620160 340720 0 0 $X=619730 $Y=340330
X490 381 472 2 3 469 NAND2X1 $T=622960 372080 1 0 $X=622530 $Y=367525
X491 381 477 2 3 476 NAND2X1 $T=625200 379920 0 0 $X=624770 $Y=379530
X564 136 8 2 3 146 AND2X1 $T=362560 387760 0 0 $X=362130 $Y=387370
X565 146 143 2 3 166 AND2X1 $T=381040 387760 1 180 $X=377250 $Y=387370
X566 166 179 2 3 176 AND2X1 $T=388880 379920 1 0 $X=388450 $Y=375365
X567 8 181 2 3 201 AND2X1 $T=411280 387760 1 180 $X=407490 $Y=387370
X568 10 214 2 3 227 AND2X1 $T=420240 340720 0 0 $X=419810 $Y=340330
X569 241 210 2 3 237 AND2X1 $T=431440 332880 1 180 $X=427650 $Y=332490
X570 242 239 2 3 214 AND2X1 $T=431440 340720 1 180 $X=427650 $Y=340330
X571 248 10 2 3 255 AND2X1 $T=434240 356400 1 0 $X=433810 $Y=351845
X572 248 253 2 3 242 AND2X1 $T=440960 356400 0 180 $X=437170 $Y=351845
X573 385 63 2 3 382 AND2X1 $T=583200 332880 0 180 $X=579410 $Y=328325
X574 401 404 2 3 394 AND2X1 $T=586560 364240 0 0 $X=586130 $Y=363850
X575 411 407 2 3 395 AND2X1 $T=593840 356400 1 180 $X=590050 $Y=356010
X576 69 387 2 3 415 AND2X1 $T=595520 332880 1 0 $X=595090 $Y=328325
X577 422 416 2 3 414 AND2X1 $T=600000 372080 1 180 $X=596210 $Y=371690
X578 436 438 2 3 441 AND2X1 $T=604480 356400 0 0 $X=604050 $Y=356010
X579 440 433 2 3 437 AND2X1 $T=606160 372080 0 0 $X=605730 $Y=371690
X580 424 451 2 3 446 AND2X1 $T=614000 340720 1 180 $X=610210 $Y=340330
X581 449 452 2 3 447 AND2X1 $T=614000 356400 1 180 $X=610210 $Y=356010
X582 443 453 2 3 448 AND2X1 $T=614000 364240 1 180 $X=610210 $Y=363850
X583 457 63 2 3 78 AND2X1 $T=616800 325040 0 0 $X=616370 $Y=324650
X584 465 459 2 3 467 AND2X1 $T=619040 348560 0 0 $X=618610 $Y=348170
X585 5 8 6 2 3 101 MUX2X1 $T=343520 426960 1 180 $X=337490 $Y=426570
X586 160 162 98 2 3 154 MUX2X1 $T=376000 340720 0 180 $X=369970 $Y=336165
X587 168 162 14 2 3 157 MUX2X1 $T=379360 356400 0 180 $X=373330 $Y=351845
X588 11 8 15 2 3 167 MUX2X1 $T=381600 403440 1 180 $X=375570 $Y=403050
X589 98 162 159 2 3 169 MUX2X1 $T=376560 332880 1 0 $X=376130 $Y=328325
X590 182 8 11 2 3 192 MUX2X1 $T=406240 411280 1 180 $X=400210 $Y=410890
X591 227 221 213 2 3 217 MUX2X1 $T=424720 332880 0 180 $X=418690 $Y=328325
X592 212 8 182 2 3 219 MUX2X1 $T=424720 411280 1 180 $X=418690 $Y=410890
X593 228 8 25 2 3 220 MUX2X1 $T=424720 419120 1 180 $X=418690 $Y=418730
X594 10 248 190 2 3 259 MUX2X1 $T=437600 364240 0 0 $X=437170 $Y=363850
X595 26 36 232 2 3 260 MUX2X1 $T=438160 325040 0 0 $X=437730 $Y=324650
X596 255 253 236 2 3 267 MUX2X1 $T=443200 356400 1 0 $X=442770 $Y=351845
X597 266 8 212 2 3 261 MUX2X1 $T=448800 403440 1 180 $X=442770 $Y=403050
X598 39 8 228 2 3 37 MUX2X1 $T=448800 419120 1 180 $X=442770 $Y=418730
X599 38 251 258 2 3 269 MUX2X1 $T=446000 325040 0 0 $X=445570 $Y=324650
X600 45 8 43 2 3 44 MUX2X1 $T=466720 426960 0 180 $X=460690 $Y=422405
X601 48 8 266 2 3 47 MUX2X1 $T=472880 395600 1 180 $X=466850 $Y=395210
X602 49 8 39 2 3 285 MUX2X1 $T=472880 419120 0 180 $X=466850 $Y=414565
X603 298 8 48 2 3 308 MUX2X1 $T=493600 395600 1 180 $X=487570 $Y=395210
X604 303 8 298 2 3 322 MUX2X1 $T=494160 395600 0 0 $X=493730 $Y=395210
X605 54 8 45 2 3 323 MUX2X1 $T=504800 419120 1 180 $X=498770 $Y=418730
X606 378 62 375 2 3 397 MUX2X1 $T=579280 403440 1 0 $X=578850 $Y=398885
X607 377 62 65 2 3 398 MUX2X1 $T=579280 419120 1 0 $X=578850 $Y=414565
X608 375 64 66 2 3 399 MUX2X1 $T=580400 426960 0 0 $X=579970 $Y=426570
X609 405 68 387 2 3 385 MUX2X1 $T=591040 332880 0 180 $X=585010 $Y=328325
X610 379 62 71 2 3 417 MUX2X1 $T=591040 395600 0 0 $X=590610 $Y=395210
X611 410 68 388 2 3 423 MUX2X1 $T=594400 356400 1 0 $X=593970 $Y=351845
X612 423 425 420 2 3 419 MUX2X1 $T=602240 340720 1 180 $X=596210 $Y=340330
X613 432 62 67 2 3 428 MUX2X1 $T=607280 395600 1 180 $X=601250 $Y=395210
X614 445 68 74 2 3 457 MUX2X1 $T=609520 325040 0 0 $X=609090 $Y=324650
X615 429 64 77 2 3 461 MUX2X1 $T=612320 419120 1 0 $X=611890 $Y=414565
X616 455 62 429 2 3 462 MUX2X1 $T=612880 403440 1 0 $X=612450 $Y=398885
X617 464 64 76 2 3 468 MUX2X1 $T=618480 419120 1 0 $X=618050 $Y=414565
X618 434 62 464 2 3 471 MUX2X1 $T=619600 403440 1 0 $X=619170 $Y=398885
X619 76 79 473 2 3 475 MUX2X1 $T=621280 426960 1 0 $X=620850 $Y=422405
X620 472 62 480 2 3 482 MUX2X1 $T=634160 379920 1 0 $X=633730 $Y=375365
X621 477 62 481 2 3 483 MUX2X1 $T=634160 387760 0 0 $X=633730 $Y=387370
X622 481 64 473 2 3 478 MUX2X1 $T=639760 411280 0 180 $X=633730 $Y=406725
X623 473 79 80 2 3 484 MUX2X1 $T=636400 419120 0 0 $X=635970 $Y=418730
X624 480 64 80 2 3 479 MUX2X1 $T=642560 411280 1 180 $X=636530 $Y=410890
X625 146 149 2 3 147 NOR2X1 $T=366480 387760 0 0 $X=366050 $Y=387370
X626 136 8 2 3 149 NOR2X1 $T=369280 387760 0 0 $X=368850 $Y=387370
X627 161 166 2 3 164 NOR2X1 $T=373200 387760 0 0 $X=372770 $Y=387370
X628 143 146 2 3 161 NOR2X1 $T=376560 379920 0 180 $X=373330 $Y=375365
X629 174 176 2 3 175 NOR2X1 $T=384960 379920 1 0 $X=384530 $Y=375365
X630 179 166 2 3 174 NOR2X1 $T=397280 379920 0 180 $X=394050 $Y=375365
X631 105 200 2 3 199 NOR2X1 $T=405680 356400 1 0 $X=405250 $Y=351845
X632 206 162 2 3 200 NOR2X1 $T=412960 356400 1 0 $X=412530 $Y=351845
X633 209 216 2 3 26 NOR2X1 $T=419680 340720 1 0 $X=419250 $Y=336165
X634 206 190 2 3 10 NOR2X1 $T=420240 364240 1 0 $X=419810 $Y=359685
X635 162 226 2 3 1 NOR2X1 $T=424160 395600 1 180 $X=420930 $Y=395210
X636 27 241 2 3 244 NOR2X1 $T=430880 332880 1 0 $X=430450 $Y=328325
X637 239 240 2 3 246 NOR2X1 $T=434240 356400 0 180 $X=431010 $Y=351845
X638 36 206 2 3 256 NOR2X1 $T=442640 340720 0 180 $X=439410 $Y=336165
X639 388 381 2 3 400 NOR2X1 $T=588800 356400 0 180 $X=585570 $Y=351845
X640 387 69 2 3 408 NOR2X1 $T=591040 332880 1 0 $X=590610 $Y=328325
X641 408 415 2 3 405 NOR2X1 $T=593840 332880 0 0 $X=593410 $Y=332490
X642 403 424 2 3 430 NOR2X1 $T=602800 340720 1 0 $X=602370 $Y=336165
X643 403 412 2 3 381 NOR2X1 $T=604480 356400 1 0 $X=604050 $Y=351845
X644 214 2 3 209 INVX2 $T=418560 340720 0 180 $X=416450 $Y=336165
X645 206 2 3 210 INVX2 $T=419120 356400 1 180 $X=417010 $Y=356010
X646 205 2 3 222 INVX2 $T=418560 387760 0 0 $X=418130 $Y=387370
X647 10 2 3 223 INVX2 $T=422480 379920 0 180 $X=420370 $Y=375365
X648 242 2 3 240 INVX2 $T=434240 356400 0 0 $X=433810 $Y=356010
X649 403 2 3 406 INVX2 $T=592160 340720 0 180 $X=590050 $Y=336165
X650 381 2 3 420 INVX2 $T=604480 356400 0 180 $X=602370 $Y=351845
X651 430 2 3 68 INVX2 $T=603360 332880 0 0 $X=602930 $Y=332490
X652 412 2 3 424 INVX2 $T=609520 340720 1 0 $X=609090 $Y=336165
X841 2 3 7 106 116 ICV_50 $T=340160 364240 0 0 $X=339730 $Y=363850
X842 2 3 114 119 117 ICV_50 $T=340160 387760 0 0 $X=339730 $Y=387370
X843 2 3 10 125 130 ICV_50 $T=350240 356400 1 0 $X=349810 $Y=351845
X844 2 3 7 103 132 ICV_50 $T=354160 340720 0 0 $X=353730 $Y=340330
X845 2 3 17 162 178 ICV_50 $T=390000 332880 1 0 $X=389570 $Y=328325
X846 2 3 16 102 196 ICV_50 $T=404560 340720 1 0 $X=404130 $Y=336165
X847 2 3 207 210 16 ICV_50 $T=411280 356400 0 0 $X=410850 $Y=356010
X848 2 3 10 221 216 ICV_50 $T=415760 340720 0 0 $X=415330 $Y=340330
X849 2 3 190 254 245 ICV_50 $T=433120 364240 0 0 $X=432690 $Y=363850
X850 2 3 251 36 241 ICV_50 $T=433680 332880 0 0 $X=433250 $Y=332490
X851 2 3 190 287 280 ICV_50 $T=467840 364240 0 0 $X=467410 $Y=363850
X852 2 3 294 296 295 ICV_50 $T=477360 340720 1 0 $X=476930 $Y=336165
X853 2 3 310 313 311 ICV_50 $T=487440 332880 0 0 $X=487010 $Y=332490
X854 2 3 7 314 294 ICV_50 $T=487440 340720 0 0 $X=487010 $Y=340330
X855 2 3 7 330 329 ICV_50 $T=500320 340720 1 0 $X=499890 $Y=336165
X856 2 3 10 340 350 ICV_50 $T=517680 403440 1 0 $X=517250 $Y=398885
X857 2 3 10 341 60 ICV_50 $T=521600 419120 0 0 $X=521170 $Y=418730
X858 2 3 412 426 422 ICV_50 $T=597760 364240 0 0 $X=597330 $Y=363850
X859 2 3 412 442 443 ICV_50 $T=606160 364240 0 0 $X=605730 $Y=363850
X895 133 135 139 2 3 134 NAND3X1 $T=353040 419120 1 0 $X=352610 $Y=414565
X896 137 142 140 2 3 141 NAND3X1 $T=363120 403440 0 180 $X=358770 $Y=398885
X897 163 13 156 2 3 12 NAND3X1 $T=375440 325040 1 180 $X=371090 $Y=324650
X898 173 13 178 2 3 177 NAND3X1 $T=384960 325040 0 0 $X=384530 $Y=324650
X899 97 171 185 2 3 184 NAND3X1 $T=392240 364240 1 0 $X=391810 $Y=359685
X900 18 13 186 2 3 19 NAND3X1 $T=392800 325040 0 0 $X=392370 $Y=324650
X901 180 13 172 2 3 183 NAND3X1 $T=396720 356400 0 180 $X=392370 $Y=351845
X902 191 13 187 2 3 188 NAND3X1 $T=401760 348560 1 180 $X=397410 $Y=348170
X903 196 13 189 2 3 193 NAND3X1 $T=404560 340720 0 180 $X=400210 $Y=336165
X904 195 13 198 2 3 24 NAND3X1 $T=403440 325040 0 0 $X=403010 $Y=324650
X905 199 13 204 2 3 3 NAND3X1 $T=408480 356400 1 0 $X=408050 $Y=351845
X906 190 206 202 2 3 208 NAND3X1 $T=415760 379920 0 180 $X=411410 $Y=375365
X907 97 225 215 2 3 224 NAND3X1 $T=423600 356400 0 180 $X=419250 $Y=351845
X908 233 10 27 2 3 225 NAND3X1 $T=427520 356400 0 180 $X=423170 $Y=351845
X909 251 221 250 2 3 249 NAND3X1 $T=438160 340720 0 180 $X=433810 $Y=336165
X910 97 264 265 2 3 263 NAND3X1 $T=443760 364240 0 0 $X=443330 $Y=363850
X911 252 268 40 2 3 270 NAND3X1 $T=448800 419120 0 0 $X=448370 $Y=418730
X912 97 273 274 2 3 275 NAND3X1 $T=462240 372080 1 180 $X=457890 $Y=371690
X913 97 278 280 2 3 277 NAND3X1 $T=462800 372080 1 0 $X=462370 $Y=367525
X914 97 279 284 2 3 46 NAND3X1 $T=463920 356400 0 0 $X=463490 $Y=356010
X915 97 276 286 2 3 281 NAND3X1 $T=464480 379920 1 0 $X=464050 $Y=375365
X916 299 309 312 2 3 315 NAND3X1 $T=489680 411280 0 0 $X=489250 $Y=410890
X917 328 318 325 2 3 326 NAND3X1 $T=504240 419120 0 180 $X=499890 $Y=414565
X918 349 321 344 2 3 347 NAND3X1 $T=520480 411280 1 180 $X=516130 $Y=410890
X919 383 63 394 2 3 389 NAND3X1 $T=579840 364240 0 0 $X=579410 $Y=363850
X920 380 63 395 2 3 393 NAND3X1 $T=580400 356400 0 0 $X=579970 $Y=356010
X921 384 392 396 2 3 386 NAND3X1 $T=580960 340720 1 0 $X=580530 $Y=336165
X922 400 63 402 2 3 3 NAND3X1 $T=589920 340720 0 0 $X=589490 $Y=340330
X923 409 63 414 2 3 413 NAND3X1 $T=591600 372080 0 0 $X=591170 $Y=371690
X924 403 424 72 2 3 421 NAND3X1 $T=602240 340720 0 180 $X=597890 $Y=336165
X925 430 427 74 2 3 396 NAND3X1 $T=604480 332880 0 180 $X=600130 $Y=328325
X926 431 63 437 2 3 435 NAND3X1 $T=602240 372080 0 0 $X=601810 $Y=371690
X927 458 63 448 2 3 460 NAND3X1 $T=614000 372080 1 0 $X=613570 $Y=367525
X928 466 63 441 2 3 463 NAND3X1 $T=621840 364240 0 180 $X=617490 $Y=359685
X929 469 63 467 2 3 474 NAND3X1 $T=628000 348560 1 180 $X=623650 $Y=348170
X930 476 63 447 2 3 470 NAND3X1 $T=628000 356400 1 180 $X=623650 $Y=356010
X972 157 153 2 3 151 OR2X1 $T=372080 348560 1 180 $X=368290 $Y=348170
X973 154 153 2 3 165 OR2X1 $T=372080 340720 0 0 $X=371650 $Y=340330
X974 169 153 2 3 170 OR2X1 $T=379360 340720 1 0 $X=378930 $Y=336165
X975 201 176 2 3 197 OR2X1 $T=407920 387760 1 180 $X=404130 $Y=387370
X976 202 176 2 3 203 OR2X1 $T=408480 379920 1 0 $X=408050 $Y=375365
X977 202 162 2 3 204 OR2X1 $T=411840 364240 0 0 $X=411410 $Y=363850
X978 210 204 2 3 215 OR2X1 $T=415760 356400 1 0 $X=415330 $Y=351845
X979 237 232 2 3 30 OR2X1 $T=430320 332880 0 180 $X=426530 $Y=328325
X980 248 206 2 3 238 OR2X1 $T=435360 348560 0 180 $X=431570 $Y=344005
X981 253 239 2 3 250 OR2X1 $T=438720 340720 1 180 $X=434930 $Y=340330
X982 256 232 2 3 258 OR2X1 $T=439280 332880 1 0 $X=438850 $Y=328325
X983 406 402 2 3 392 OR2X1 $T=589920 340720 1 180 $X=586130 $Y=340330
X984 70 387 2 3 418 OR2X1 $T=593840 325040 0 0 $X=593410 $Y=324650
X985 72 412 2 3 402 OR2X1 $T=598320 340720 0 180 $X=594530 $Y=336165
X986 73 418 2 3 427 OR2X1 $T=598880 325040 0 0 $X=598450 $Y=324650
X987 446 425 2 3 456 OR2X1 $T=617360 340720 1 180 $X=613570 $Y=340330
X988 162 2 3 190 INVX8 $T=423600 379920 1 0 $X=423170 $Y=375365
X989 229 2 3 7 INVX8 $T=427520 387760 1 0 $X=427090 $Y=383205
X990 2 72 ANTENNA $T=596640 332880 0 0 $X=596210 $Y=332490
X991 2 72 ANTENNA $T=597760 332880 0 0 $X=597330 $Y=332490
X992 430 73 3 2 75 XOR2X1 $T=602240 325040 0 0 $X=601810 $Y=324650
X993 415 74 3 2 445 XOR2X1 $T=606720 332880 1 0 $X=606290 $Y=328325
.ENDS
***************************************
.SUBCKT ICV_46
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT INVX1 A VSS VDD Z
** N=6 EP=4 IP=0 FDC=2
M0 Z A VSS VSS N L=1.8e-07 W=2.2e-07 $X=740 $Y=760 $D=0
M1 Z A VDD VDD P L=1.8e-07 W=4.4e-07 $X=740 $Y=2715 $D=16
.ENDS
***************************************
.SUBCKT ICV_47 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111
** N=383 EP=111 IP=4039 FDC=4662
X32 123 105 106 2 1 2 121 DFFQSRX1 $T=314400 458320 1 0 $X=313970 $Y=453765
X33 120 105 106 2 1 2 122 DFFQSRX1 $T=314400 474000 0 0 $X=313970 $Y=473610
X34 117 105 106 2 1 2 3 DFFQSRX1 $T=349120 497520 0 180 $X=323490 $Y=492965
X35 124 105 106 2 1 2 4 DFFQSRX1 $T=353040 442640 0 180 $X=327410 $Y=438085
X36 118 105 106 2 1 2 5 DFFQSRX1 $T=353600 434800 1 180 $X=327970 $Y=434410
X37 119 105 106 2 1 2 114 DFFQSRX1 $T=353600 458320 1 180 $X=327970 $Y=457930
X38 125 105 106 2 1 2 115 DFFQSRX1 $T=353600 466160 0 180 $X=327970 $Y=461605
X39 126 105 106 2 1 2 116 DFFQSRX1 $T=353600 489680 1 180 $X=327970 $Y=489290
X40 162 105 106 2 1 2 137 DFFQSRX1 $T=345200 481840 1 0 $X=344770 $Y=477285
X41 130 105 106 2 1 2 129 DFFQSRX1 $T=345200 481840 0 0 $X=344770 $Y=481450
X42 128 105 106 2 1 2 132 DFFQSRX1 $T=353600 434800 0 0 $X=353170 $Y=434410
X43 141 105 106 2 1 2 127 DFFQSRX1 $T=380480 466160 0 180 $X=354850 $Y=461605
X44 139 105 106 2 1 2 131 DFFQSRX1 $T=386640 442640 0 180 $X=361010 $Y=438085
X45 150 105 106 2 1 2 133 DFFQSRX1 $T=386640 458320 1 180 $X=361010 $Y=457930
X46 154 105 106 2 1 2 134 DFFQSRX1 $T=386640 489680 1 180 $X=361010 $Y=489290
X47 140 105 106 2 1 2 135 DFFQSRX1 $T=386640 497520 0 180 $X=361010 $Y=492965
X48 159 105 106 2 1 2 138 DFFQSRX1 $T=397280 481840 0 180 $X=371650 $Y=477285
X49 231 105 106 2 1 2 144 DFFQSRX1 $T=400640 481840 1 180 $X=375010 $Y=481450
X50 168 105 106 2 1 2 157 DFFQSRX1 $T=380480 466160 1 0 $X=380050 $Y=461605
X51 164 105 106 2 1 2 163 DFFQSRX1 $T=381600 434800 0 0 $X=381170 $Y=434410
X52 169 105 106 2 1 2 160 DFFQSRX1 $T=416320 442640 0 180 $X=390690 $Y=438085
X53 218 105 106 2 1 2 161 DFFQSRX1 $T=416880 489680 1 180 $X=391250 $Y=489290
X54 173 105 106 2 1 2 177 DFFQSRX1 $T=402320 481840 0 0 $X=401890 $Y=481450
X55 194 105 106 2 1 2 170 DFFQSRX1 $T=428080 481840 0 180 $X=402450 $Y=477285
X56 175 105 106 2 1 2 184 DFFQSRX1 $T=406240 458320 0 0 $X=405810 $Y=457930
X57 183 105 106 2 1 2 180 DFFQSRX1 $T=406240 466160 1 0 $X=405810 $Y=461605
X58 179 105 106 2 1 2 38 DFFQSRX1 $T=406240 497520 1 0 $X=405810 $Y=492965
X59 188 105 106 2 1 2 193 DFFQSRX1 $T=408480 434800 0 0 $X=408050 $Y=434410
X60 192 105 106 2 1 2 185 DFFQSRX1 $T=442080 489680 1 180 $X=416450 $Y=489290
X61 206 105 106 2 1 2 191 DFFQSRX1 $T=447120 442640 0 180 $X=421490 $Y=438085
X62 204 105 106 2 1 2 209 DFFQSRX1 $T=433120 481840 0 0 $X=432690 $Y=481450
X63 226 105 106 2 1 2 52 DFFQSRX1 $T=436480 481840 1 0 $X=436050 $Y=477285
X64 202 105 106 2 1 2 197 DFFQSRX1 $T=437040 458320 0 0 $X=436610 $Y=457930
X65 216 105 106 2 1 2 211 DFFQSRX1 $T=437040 497520 1 0 $X=436610 $Y=492965
X66 108 105 106 2 1 2 45 DFFQSRX1 $T=472320 442640 0 180 $X=446690 $Y=438085
X67 229 105 106 2 1 2 214 DFFQSRX1 $T=472880 466160 0 180 $X=447250 $Y=461605
X68 219 105 106 2 1 2 217 DFFQSRX1 $T=475120 489680 1 180 $X=449490 $Y=489290
X69 109 105 106 2 1 2 48 DFFQSRX1 $T=477360 434800 1 180 $X=451730 $Y=434410
X70 107 105 106 2 1 2 63 DFFQSRX1 $T=463360 481840 0 0 $X=462930 $Y=481450
X71 247 105 106 2 1 2 254 DFFQSRX1 $T=466720 481840 1 0 $X=466290 $Y=477285
X72 245 105 106 2 1 2 251 DFFQSRX1 $T=472880 458320 0 0 $X=472450 $Y=457930
X73 253 105 106 2 1 2 252 DFFQSRX1 $T=472880 466160 1 0 $X=472450 $Y=461605
X74 255 105 106 2 1 2 238 DFFQSRX1 $T=502560 434800 1 180 $X=476930 $Y=434410
X75 262 105 106 2 1 2 246 DFFQSRX1 $T=508160 442640 0 180 $X=482530 $Y=438085
X76 264 105 106 2 1 2 248 DFFQSRX1 $T=508160 489680 1 180 $X=482530 $Y=489290
X77 260 105 106 2 1 2 60 DFFQSRX1 $T=508160 497520 0 180 $X=482530 $Y=492965
X78 223 105 106 2 1 2 227 DFFQSRX1 $T=493600 481840 1 0 $X=493170 $Y=477285
X79 259 105 106 2 1 2 261 DFFQSRX1 $T=493600 481840 0 0 $X=493170 $Y=481450
X80 270 105 106 2 1 2 258 DFFQSRX1 $T=498080 458320 0 0 $X=497650 $Y=457930
X81 110 105 106 2 1 2 66 DFFQSRX1 $T=502560 434800 0 0 $X=502130 $Y=434410
X82 286 105 106 2 1 2 276 DFFQSRX1 $T=536720 489680 1 180 $X=511090 $Y=489290
X83 293 105 106 2 1 2 277 DFFQSRX1 $T=537280 466160 0 180 $X=511650 $Y=461605
X84 281 105 106 2 1 2 273 DFFQSRX1 $T=537280 497520 0 180 $X=511650 $Y=492965
X85 282 105 106 2 1 2 70 DFFQSRX1 $T=538400 442640 0 180 $X=512770 $Y=438085
X86 266 105 106 2 1 2 279 DFFQSRX1 $T=524400 481840 1 0 $X=523970 $Y=477285
X87 295 105 106 2 1 2 76 DFFQSRX1 $T=549600 481840 1 180 $X=523970 $Y=481450
X88 291 105 106 2 1 2 79 DFFQSRX1 $T=528320 434800 0 0 $X=527890 $Y=434410
X89 235 105 106 2 1 2 241 DFFQSRX1 $T=528320 458320 0 0 $X=527890 $Y=457930
X90 236 105 106 2 1 2 56 DFFQSRX1 $T=561920 489680 1 180 $X=536290 $Y=489290
X91 111 105 106 2 1 2 81 DFFQSRX1 $T=562480 497520 0 180 $X=536850 $Y=492965
X92 240 105 106 2 1 2 244 DFFQSRX1 $T=561920 489680 0 0 $X=561490 $Y=489290
X93 54 105 106 2 1 2 233 DFFQSRX1 $T=562480 497520 1 0 $X=562050 $Y=492965
X94 301 105 106 2 1 2 82 DFFQSRX1 $T=592720 458320 1 180 $X=567090 $Y=457930
X95 312 105 106 2 1 2 296 DFFQSRX1 $T=592720 466160 0 180 $X=567090 $Y=461605
X96 307 105 106 2 1 2 297 DFFQSRX1 $T=593840 442640 0 180 $X=568210 $Y=438085
X97 310 105 106 2 1 2 83 DFFQSRX1 $T=594400 434800 1 180 $X=568770 $Y=434410
X98 348 105 106 2 1 2 318 DFFQSRX1 $T=613440 481840 1 180 $X=587810 $Y=481450
X99 321 105 106 2 1 2 89 DFFQSRX1 $T=592720 458320 0 0 $X=592290 $Y=457930
X100 335 105 106 2 1 2 327 DFFQSRX1 $T=592720 466160 1 0 $X=592290 $Y=461605
X101 333 105 106 2 1 2 320 DFFQSRX1 $T=593840 442640 1 0 $X=593410 $Y=438085
X102 346 105 106 2 1 2 329 DFFQSRX1 $T=625200 489680 1 180 $X=599570 $Y=489290
X103 349 105 106 2 1 2 96 DFFQSRX1 $T=625200 497520 0 180 $X=599570 $Y=492965
X104 347 105 106 2 1 2 330 DFFQSRX1 $T=626320 434800 1 180 $X=600690 $Y=434410
X105 350 105 106 2 1 2 101 DFFQSRX1 $T=619600 442640 1 0 $X=619170 $Y=438085
X106 356 105 106 2 1 2 103 DFFQSRX1 $T=627440 434800 0 0 $X=627010 $Y=434410
X107 359 105 106 2 1 2 351 DFFQSRX1 $T=652640 442640 1 180 $X=627010 $Y=442250
X108 360 105 106 2 1 2 358 DFFQSRX1 $T=628560 458320 1 0 $X=628130 $Y=453765
X109 362 105 106 2 1 2 352 DFFQSRX1 $T=653760 466160 0 180 $X=628130 $Y=461605
X110 357 105 106 2 1 2 361 DFFQSRX1 $T=629120 474000 0 0 $X=628690 $Y=473610
X111 363 105 106 2 1 2 353 DFFQSRX1 $T=654320 481840 0 180 $X=628690 $Y=477285
X112 364 105 106 2 1 2 354 DFFQSRX1 $T=654320 489680 0 180 $X=628690 $Y=485125
X113 365 105 106 2 1 2 355 DFFQSRX1 $T=654320 497520 0 180 $X=628690 $Y=492965
X253 14 13 1 2 136 NAND2X1 $T=370400 434800 0 180 $X=367170 $Y=430245
X254 18 138 1 2 143 NAND2X1 $T=377120 458320 0 180 $X=373890 $Y=453765
X255 14 133 1 2 146 NAND2X1 $T=381600 434800 1 180 $X=378370 $Y=434410
X256 18 133 1 2 145 NAND2X1 $T=383280 458320 0 180 $X=380050 $Y=453765
X257 14 138 1 2 153 NAND2X1 $T=386080 474000 0 180 $X=382850 $Y=469445
X258 25 132 1 2 142 NAND2X1 $T=388320 434800 0 180 $X=385090 $Y=430245
X259 25 131 1 2 155 NAND2X1 $T=386080 442640 0 0 $X=385650 $Y=442250
X260 18 26 1 2 151 NAND2X1 $T=389440 442640 0 180 $X=386210 $Y=438085
X261 18 157 1 2 156 NAND2X1 $T=386640 458320 0 0 $X=386210 $Y=457930
X262 25 135 1 2 147 NAND2X1 $T=387200 497520 1 0 $X=386770 $Y=492965
X263 25 20 1 2 148 NAND2X1 $T=388880 442640 0 0 $X=388450 $Y=442250
X264 25 127 1 2 158 NAND2X1 $T=390000 497520 1 0 $X=389570 $Y=492965
X265 18 163 1 2 149 NAND2X1 $T=390560 434800 1 0 $X=390130 $Y=430245
X266 25 28 1 2 152 NAND2X1 $T=393360 434800 1 0 $X=392930 $Y=430245
X267 14 157 1 2 165 NAND2X1 $T=393360 458320 0 0 $X=392930 $Y=457930
X268 14 163 1 2 167 NAND2X1 $T=393920 450480 1 0 $X=393490 $Y=445925
X269 25 134 1 2 166 NAND2X1 $T=397840 489680 1 0 $X=397410 $Y=485125
X270 25 137 1 2 171 NAND2X1 $T=404560 489680 1 0 $X=404130 $Y=485125
X271 25 160 1 2 172 NAND2X1 $T=405120 442640 0 0 $X=404690 $Y=442250
X272 14 180 1 2 181 NAND2X1 $T=414640 458320 0 180 $X=411410 $Y=453765
X273 18 180 1 2 178 NAND2X1 $T=416880 489680 0 180 $X=413650 $Y=485125
X274 25 31 1 2 182 NAND2X1 $T=414640 434800 1 0 $X=414210 $Y=430245
X275 14 184 1 2 176 NAND2X1 $T=414640 450480 1 0 $X=414210 $Y=445925
X276 18 170 1 2 174 NAND2X1 $T=420800 474000 0 180 $X=417570 $Y=469445
X277 14 170 1 2 189 NAND2X1 $T=421920 489680 0 180 $X=418690 $Y=485125
X278 18 184 1 2 187 NAND2X1 $T=420240 442640 0 0 $X=419810 $Y=442250
X279 18 193 1 2 186 NAND2X1 $T=420240 450480 1 0 $X=419810 $Y=445925
X280 14 193 1 2 190 NAND2X1 $T=428080 434800 0 180 $X=424850 $Y=430245
X281 14 36 1 2 195 NAND2X1 $T=428080 505360 1 0 $X=427650 $Y=500805
X282 14 197 1 2 198 NAND2X1 $T=433120 450480 0 180 $X=429890 $Y=445925
X283 25 177 1 2 196 NAND2X1 $T=430880 489680 1 0 $X=430450 $Y=485125
X284 14 39 1 2 199 NAND2X1 $T=434240 434800 0 180 $X=431010 $Y=430245
X285 25 185 1 2 200 NAND2X1 $T=431440 497520 1 0 $X=431010 $Y=492965
X286 18 197 1 2 201 NAND2X1 $T=434800 474000 0 180 $X=431570 $Y=469445
X287 18 39 1 2 203 NAND2X1 $T=436480 434800 1 180 $X=433250 $Y=434410
X288 25 33 1 2 207 NAND2X1 $T=438160 442640 0 0 $X=437730 $Y=442250
X289 18 211 1 2 205 NAND2X1 $T=440400 474000 1 0 $X=439970 $Y=469445
X290 14 191 1 2 208 NAND2X1 $T=442640 450480 1 0 $X=442210 $Y=445925
X291 14 211 1 2 212 NAND2X1 $T=446000 489680 1 180 $X=442770 $Y=489290
X292 18 191 1 2 210 NAND2X1 $T=447120 434800 0 180 $X=443890 $Y=430245
X293 18 44 1 2 213 NAND2X1 $T=447680 442640 1 180 $X=444450 $Y=442250
X294 18 214 1 2 46 NAND2X1 $T=447120 434800 0 0 $X=446690 $Y=434410
X295 14 144 1 2 220 NAND2X1 $T=453840 489680 1 0 $X=453410 $Y=485125
X296 14 214 1 2 222 NAND2X1 $T=457200 450480 0 180 $X=453970 $Y=445925
X297 18 217 1 2 221 NAND2X1 $T=454400 466160 0 0 $X=453970 $Y=465770
X298 25 209 1 2 215 NAND2X1 $T=460560 497520 1 180 $X=457330 $Y=497130
X299 25 161 1 2 225 NAND2X1 $T=462800 505360 0 180 $X=459570 $Y=500805
X300 14 217 1 2 224 NAND2X1 $T=460560 442640 0 0 $X=460130 $Y=442250
X301 18 144 1 2 228 NAND2X1 $T=463360 466160 1 180 $X=460130 $Y=465770
X302 14 56 1 2 232 NAND2X1 $T=464480 497520 0 0 $X=464050 $Y=497130
X303 25 227 1 2 230 NAND2X1 $T=467280 489680 1 0 $X=466850 $Y=485125
X304 25 233 1 2 234 NAND2X1 $T=474000 505360 1 0 $X=473570 $Y=500805
X305 25 241 1 2 239 NAND2X1 $T=476240 474000 1 0 $X=475810 $Y=469445
X306 14 251 1 2 249 NAND2X1 $T=482960 442640 0 0 $X=482530 $Y=442250
X307 18 252 1 2 243 NAND2X1 $T=484080 458320 1 0 $X=483650 $Y=453765
X308 14 252 1 2 250 NAND2X1 $T=489680 458320 0 180 $X=486450 $Y=453765
X309 18 251 1 2 237 NAND2X1 $T=488560 489680 1 0 $X=488130 $Y=485125
X310 25 244 1 2 256 NAND2X1 $T=493600 481840 1 180 $X=490370 $Y=481450
X311 18 258 1 2 257 NAND2X1 $T=491360 489680 1 0 $X=490930 $Y=485125
X312 25 66 1 2 242 NAND2X1 $T=495280 434800 1 0 $X=494850 $Y=430245
X313 25 254 1 2 263 NAND2X1 $T=500320 474000 0 180 $X=497090 $Y=469445
X314 14 258 1 2 267 NAND2X1 $T=505920 450480 1 180 $X=502690 $Y=450090
X315 18 67 1 2 265 NAND2X1 $T=503680 505360 1 0 $X=503250 $Y=500805
X316 25 238 1 2 269 NAND2X1 $T=509280 434800 0 180 $X=506050 $Y=430245
X317 25 246 1 2 271 NAND2X1 $T=508160 442640 1 0 $X=507730 $Y=438085
X318 25 273 1 2 272 NAND2X1 $T=508160 489680 0 0 $X=507730 $Y=489290
X319 25 69 1 2 275 NAND2X1 $T=512080 434800 0 180 $X=508850 $Y=430245
X320 25 248 1 2 274 NAND2X1 $T=509280 497520 1 0 $X=508850 $Y=492965
X321 14 279 1 2 268 NAND2X1 $T=510400 474000 1 0 $X=509970 $Y=469445
X322 25 261 1 2 278 NAND2X1 $T=510960 505360 1 0 $X=510530 $Y=500805
X323 18 279 1 2 284 NAND2X1 $T=516000 458320 1 0 $X=515570 $Y=453765
X324 18 277 1 2 283 NAND2X1 $T=518800 466160 1 180 $X=515570 $Y=465770
X325 14 277 1 2 285 NAND2X1 $T=516560 450480 1 0 $X=516130 $Y=445925
X326 14 70 1 2 280 NAND2X1 $T=520480 442640 1 180 $X=517250 $Y=442250
X327 14 276 1 2 288 NAND2X1 $T=521600 481840 0 0 $X=521170 $Y=481450
X328 14 76 1 2 290 NAND2X1 $T=521600 489680 1 0 $X=521170 $Y=485125
X329 18 276 1 2 292 NAND2X1 $T=522720 466160 0 0 $X=522290 $Y=465770
X330 18 78 1 2 294 NAND2X1 $T=523280 458320 0 0 $X=522850 $Y=457930
X331 14 79 1 2 289 NAND2X1 $T=524960 434800 1 0 $X=524530 $Y=430245
X332 14 80 1 2 287 NAND2X1 $T=524960 505360 1 0 $X=524530 $Y=500805
X333 303 299 1 2 301 NAND2X1 $T=577600 474000 1 180 $X=574370 $Y=473610
X334 304 87 1 2 302 NAND2X1 $T=577600 505360 0 180 $X=574370 $Y=500805
X335 84 305 1 2 300 NAND2X1 $T=575920 489680 1 0 $X=575490 $Y=485125
X336 304 82 1 2 303 NAND2X1 $T=579280 481840 1 0 $X=578850 $Y=477285
X337 85 84 1 2 308 NAND2X1 $T=580400 505360 1 0 $X=579970 $Y=500805
X338 306 305 1 2 304 NAND2X1 $T=582080 489680 1 0 $X=581650 $Y=485125
X339 313 311 1 2 312 NAND2X1 $T=587120 474000 1 180 $X=583890 $Y=473610
X340 90 315 1 2 311 NAND2X1 $T=584880 481840 1 0 $X=584450 $Y=477285
X341 302 308 1 2 91 NAND2X1 $T=588240 505360 0 180 $X=585010 $Y=500805
X342 91 296 1 2 313 NAND2X1 $T=592720 481840 0 180 $X=589490 $Y=477285
X343 322 324 1 2 314 NAND2X1 $T=592720 481840 1 0 $X=592290 $Y=477285
X344 96 318 1 2 324 NAND2X1 $T=593840 497520 1 0 $X=593410 $Y=492965
X345 327 329 1 2 328 NAND2X1 $T=597200 474000 1 0 $X=596770 $Y=469445
X346 334 337 1 2 335 NAND2X1 $T=603360 474000 0 0 $X=602930 $Y=473610
X347 325 327 1 2 336 NAND2X1 $T=603360 489680 1 0 $X=602930 $Y=485125
X348 91 327 1 2 334 NAND2X1 $T=606720 481840 1 0 $X=606290 $Y=477285
X349 90 338 1 2 340 NAND2X1 $T=610080 505360 0 180 $X=606850 $Y=500805
X350 91 318 1 2 341 NAND2X1 $T=611760 497520 1 180 $X=608530 $Y=497130
X351 91 329 1 2 343 NAND2X1 $T=610080 474000 0 0 $X=609650 $Y=473610
X352 91 96 1 2 344 NAND2X1 $T=613440 505360 0 180 $X=610210 $Y=500805
X353 345 343 1 2 346 NAND2X1 $T=615680 474000 1 180 $X=612450 $Y=473610
X354 341 339 1 2 348 NAND2X1 $T=616240 497520 1 180 $X=613010 $Y=497130
X355 344 340 1 2 349 NAND2X1 $T=616240 505360 0 180 $X=613010 $Y=500805
X448 3 7 6 1 2 117 MUX2X1 $T=334560 505360 0 180 $X=328530 $Y=500805
X449 5 9 114 1 2 118 MUX2X1 $T=343520 434800 0 180 $X=337490 $Y=430245
X450 122 8 114 1 2 119 MUX2X1 $T=344080 442640 1 180 $X=338050 $Y=442250
X451 115 8 4 1 2 124 MUX2X1 $T=338480 450480 1 0 $X=338050 $Y=445925
X452 122 7 116 1 2 120 MUX2X1 $T=344080 466160 1 180 $X=338050 $Y=465770
X453 115 7 122 1 2 125 MUX2X1 $T=338480 474000 1 0 $X=338050 $Y=469445
X454 116 7 10 1 2 126 MUX2X1 $T=339040 489680 1 0 $X=338610 $Y=485125
X455 116 8 121 1 2 123 MUX2X1 $T=345200 458320 0 180 $X=339170 $Y=453765
X456 10 7 11 1 2 12 MUX2X1 $T=352480 497520 0 0 $X=352050 $Y=497130
X457 10 8 129 1 2 130 MUX2X1 $T=354160 489680 0 0 $X=353730 $Y=489290
X458 132 9 121 1 2 128 MUX2X1 $T=363120 442640 1 180 $X=357090 $Y=442250
X459 131 9 132 1 2 139 MUX2X1 $T=378240 442640 1 180 $X=372210 $Y=442250
X460 135 9 15 1 2 140 MUX2X1 $T=378240 497520 1 180 $X=372210 $Y=497130
X461 127 9 129 1 2 141 MUX2X1 $T=378800 489680 0 180 $X=372770 $Y=485125
X462 20 9 19 1 2 17 MUX2X1 $T=381600 434800 0 180 $X=375570 $Y=430245
X463 134 9 127 1 2 154 MUX2X1 $T=392240 489680 0 180 $X=386210 $Y=485125
X464 137 9 135 1 2 162 MUX2X1 $T=397840 489680 0 180 $X=391810 $Y=485125
X465 160 9 131 1 2 169 MUX2X1 $T=402880 434800 0 180 $X=396850 $Y=430245
X466 31 9 20 1 2 30 MUX2X1 $T=408480 434800 0 180 $X=402450 $Y=430245
X467 177 9 134 1 2 173 MUX2X1 $T=413520 489680 0 180 $X=407490 $Y=485125
X468 33 9 160 1 2 32 MUX2X1 $T=414080 434800 0 180 $X=408050 $Y=430245
X469 185 9 137 1 2 192 MUX2X1 $T=427520 489680 0 180 $X=421490 $Y=485125
X470 209 9 177 1 2 204 MUX2X1 $T=440960 489680 0 180 $X=434930 $Y=485125
X471 161 9 185 1 2 218 MUX2X1 $T=456080 505360 0 180 $X=450050 $Y=500805
X472 227 9 209 1 2 223 MUX2X1 $T=462240 489680 0 180 $X=456210 $Y=485125
X473 52 9 33 1 2 226 MUX2X1 $T=465040 434800 0 180 $X=459010 $Y=430245
X474 233 9 161 1 2 54 MUX2X1 $T=470080 505360 0 180 $X=464050 $Y=500805
X475 241 9 227 1 2 235 MUX2X1 $T=481280 489680 0 180 $X=475250 $Y=485125
X476 244 9 233 1 2 240 MUX2X1 $T=483520 497520 1 180 $X=477490 $Y=497130
X477 254 9 241 1 2 247 MUX2X1 $T=488560 489680 0 180 $X=482530 $Y=485125
X478 238 9 64 1 2 255 MUX2X1 $T=494160 434800 0 180 $X=488130 $Y=430245
X479 261 9 244 1 2 259 MUX2X1 $T=499760 489680 0 180 $X=493730 $Y=485125
X480 246 9 238 1 2 262 MUX2X1 $T=504240 434800 0 180 $X=498210 $Y=430245
X481 248 9 254 1 2 264 MUX2X1 $T=505360 489680 0 180 $X=499330 $Y=485125
X482 273 9 261 1 2 281 MUX2X1 $T=510400 489680 1 0 $X=509970 $Y=485125
X483 71 9 69 1 2 73 MUX2X1 $T=513200 434800 1 0 $X=512770 $Y=430245
X484 83 88 297 1 2 310 MUX2X1 $T=579840 434800 1 0 $X=579410 $Y=430245
X485 297 90 89 1 2 307 MUX2X1 $T=585440 442640 1 180 $X=579410 $Y=442250
X486 89 90 320 1 2 321 MUX2X1 $T=588240 442640 0 0 $X=587810 $Y=442250
X487 93 88 320 1 2 97 MUX2X1 $T=591040 434800 1 0 $X=590610 $Y=430245
X488 320 90 330 1 2 333 MUX2X1 $T=598880 442640 0 0 $X=598450 $Y=442250
X489 99 88 330 1 2 100 MUX2X1 $T=601680 434800 1 0 $X=601250 $Y=430245
X490 330 90 101 1 2 347 MUX2X1 $T=609520 434800 1 0 $X=609090 $Y=430245
X491 101 90 102 1 2 350 MUX2X1 $T=615120 434800 1 0 $X=614690 $Y=430245
X492 351 90 358 1 2 359 MUX2X1 $T=636400 450480 0 0 $X=635970 $Y=450090
X493 103 90 351 1 2 356 MUX2X1 $T=642560 434800 0 180 $X=636530 $Y=430245
X494 352 90 361 1 2 362 MUX2X1 $T=639200 466160 0 0 $X=638770 $Y=465770
X495 361 90 353 1 2 357 MUX2X1 $T=644800 474000 0 180 $X=638770 $Y=469445
X496 353 90 354 1 2 363 MUX2X1 $T=639200 481840 0 0 $X=638770 $Y=481450
X497 354 90 355 1 2 364 MUX2X1 $T=639200 489680 0 0 $X=638770 $Y=489290
X498 355 90 104 1 2 365 MUX2X1 $T=639200 505360 1 0 $X=638770 $Y=500805
X499 358 90 352 1 2 360 MUX2X1 $T=647600 450480 1 180 $X=641570 $Y=450090
X500 314 317 1 2 88 NOR2X1 $T=585440 481840 0 0 $X=585010 $Y=481450
X501 95 324 1 2 325 NOR2X1 $T=597200 489680 1 180 $X=593970 $Y=489290
X502 328 326 1 2 323 NOR2X1 $T=598880 474000 1 180 $X=595650 $Y=473610
X503 329 327 1 2 322 NOR2X1 $T=600560 489680 0 180 $X=597330 $Y=485125
X504 85 1 2 305 INVX2 $T=577600 497520 0 0 $X=577170 $Y=497130
X505 318 1 2 92 INVX2 $T=600000 505360 0 180 $X=597890 $Y=500805
X506 325 1 2 326 INVX2 $T=602240 489680 0 180 $X=600130 $Y=485125
X645 136 142 143 1 2 16 NAND3X1 $T=372080 434800 1 0 $X=371650 $Y=430245
X646 146 148 151 1 2 150 NAND3X1 $T=379360 442640 0 0 $X=378930 $Y=442250
X647 23 147 145 1 2 21 NAND3X1 $T=383280 489680 0 180 $X=378930 $Y=485125
X648 24 152 149 1 2 22 NAND3X1 $T=385520 434800 0 180 $X=381170 $Y=430245
X649 153 158 27 1 2 159 NAND3X1 $T=386640 489680 0 0 $X=386210 $Y=489290
X650 167 155 156 1 2 164 NAND3X1 $T=396720 450480 1 180 $X=392370 $Y=450090
X651 165 166 29 1 2 168 NAND3X1 $T=393360 474000 1 0 $X=392930 $Y=469445
X652 176 172 174 1 2 175 NAND3X1 $T=412960 450480 0 180 $X=408610 $Y=445925
X653 34 171 178 1 2 179 NAND3X1 $T=415760 497520 1 180 $X=411410 $Y=497130
X654 181 182 186 1 2 183 NAND3X1 $T=414640 458320 1 0 $X=414210 $Y=453765
X655 190 35 187 1 2 188 NAND3X1 $T=423040 434800 0 180 $X=418690 $Y=430245
X656 189 196 37 1 2 194 NAND3X1 $T=427520 481840 0 0 $X=427090 $Y=481450
X657 198 40 203 1 2 202 NAND3X1 $T=430880 442640 0 0 $X=430450 $Y=442250
X658 195 200 201 1 2 41 NAND3X1 $T=430880 505360 1 0 $X=430450 $Y=500805
X659 199 42 210 1 2 43 NAND3X1 $T=436480 434800 0 0 $X=436050 $Y=434410
X660 208 207 205 1 2 206 NAND3X1 $T=440400 450480 0 180 $X=436050 $Y=445925
X661 212 215 47 1 2 216 NAND3X1 $T=446000 489680 0 0 $X=445570 $Y=489290
X662 224 49 213 1 2 219 NAND3X1 $T=458320 442640 1 180 $X=453970 $Y=442250
X663 51 225 221 1 2 50 NAND3X1 $T=460000 505360 0 180 $X=455650 $Y=500805
X664 222 53 228 1 2 229 NAND3X1 $T=460000 450480 1 0 $X=459570 $Y=445925
X665 220 230 55 1 2 231 NAND3X1 $T=462240 489680 1 0 $X=461810 $Y=485125
X666 232 234 237 1 2 236 NAND3X1 $T=473440 497520 0 0 $X=473010 $Y=497130
X667 57 242 243 1 2 58 NAND3X1 $T=477920 434800 1 0 $X=477490 $Y=430245
X668 249 61 59 1 2 245 NAND3X1 $T=485760 434800 0 180 $X=481410 $Y=430245
X669 250 239 62 1 2 253 NAND3X1 $T=484080 474000 1 0 $X=483650 $Y=469445
X670 65 256 257 1 2 260 NAND3X1 $T=494720 497520 0 0 $X=494290 $Y=497130
X671 268 263 265 1 2 266 NAND3X1 $T=507600 474000 1 180 $X=503250 $Y=473610
X672 267 269 68 1 2 270 NAND3X1 $T=505920 450480 1 0 $X=505490 $Y=445925
X673 280 275 284 1 2 282 NAND3X1 $T=513760 442640 0 0 $X=513330 $Y=442250
X674 287 278 283 1 2 74 NAND3X1 $T=520480 505360 0 180 $X=516130 $Y=500805
X675 288 274 72 1 2 286 NAND3X1 $T=521600 489680 0 180 $X=517250 $Y=485125
X676 289 75 292 1 2 291 NAND3X1 $T=521040 434800 1 0 $X=520610 $Y=430245
X677 285 271 77 1 2 293 NAND3X1 $T=521600 450480 1 0 $X=521170 $Y=445925
X678 290 272 294 1 2 295 NAND3X1 $T=524400 489680 1 0 $X=523970 $Y=485125
X679 2 298 300 1 2 1 NAND3X1 $T=572000 489680 1 0 $X=571570 $Y=485125
X680 84 85 86 1 2 299 NAND3X1 $T=572000 497520 0 0 $X=571570 $Y=497130
X681 304 308 86 1 2 309 NAND3X1 $T=585440 497520 1 180 $X=581090 $Y=497130
X682 319 305 296 1 2 316 NAND3X1 $T=591600 489680 1 180 $X=587250 $Y=489290
X683 95 94 92 1 2 319 NAND3X1 $T=594960 505360 0 180 $X=590610 $Y=500805
X684 86 306 1 2 298 OR2X1 $T=582080 489680 0 180 $X=578290 $Y=485125
X685 306 316 1 2 317 OR2X1 $T=585440 489680 1 0 $X=585010 $Y=485125
X686 331 309 1 2 337 OR2X1 $T=603360 481840 1 0 $X=602930 $Y=477285
X687 332 309 1 2 339 OR2X1 $T=603920 497520 0 0 $X=603490 $Y=497130
X688 309 342 1 2 345 OR2X1 $T=609520 481840 1 0 $X=609090 $Y=477285
X689 309 1 2 90 INVX8 $T=587680 497520 0 0 $X=587250 $Y=497130
X690 323 296 2 1 315 XOR2X1 $T=594400 474000 1 180 $X=587810 $Y=473610
X691 326 327 2 1 331 XOR2X1 $T=596080 481840 1 0 $X=595650 $Y=477285
X692 95 318 2 1 332 XOR2X1 $T=597200 497520 0 0 $X=596770 $Y=497130
X693 98 96 2 1 338 XOR2X1 $T=600000 505360 1 0 $X=599570 $Y=500805
X694 336 329 2 1 342 XOR2X1 $T=607840 489680 1 0 $X=607410 $Y=485125
X725 84 1 2 306 INVX1 $T=578160 481840 0 0 $X=577730 $Y=481450
.ENDS
***************************************
.SUBCKT ICV_39
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_45 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 54
** N=374 EP=53 IP=4449 FDC=5598
X43 149 47 48 2 1 2 56 DFFQSRX1 $T=339600 513200 0 180 $X=313970 $Y=508645
X44 143 47 48 2 1 2 72 DFFQSRX1 $T=314400 528880 1 0 $X=313970 $Y=524325
X45 64 47 48 2 1 2 73 DFFQSRX1 $T=314400 536720 0 0 $X=313970 $Y=536330
X46 79 47 48 2 1 2 57 DFFQSRX1 $T=339600 544560 0 180 $X=313970 $Y=540005
X47 65 47 48 2 1 2 68 DFFQSRX1 $T=314400 552400 0 0 $X=313970 $Y=552010
X48 220 47 48 2 1 2 58 DFFQSRX1 $T=339600 560240 0 180 $X=313970 $Y=555685
X49 66 47 48 2 1 2 69 DFFQSRX1 $T=314400 560240 0 0 $X=313970 $Y=559850
X50 209 47 48 2 1 2 74 DFFQSRX1 $T=314400 583760 0 0 $X=313970 $Y=583370
X51 70 47 48 2 1 2 75 DFFQSRX1 $T=314400 591600 0 0 $X=313970 $Y=591210
X52 104 47 48 2 1 2 59 DFFQSRX1 $T=339600 599440 0 180 $X=313970 $Y=594885
X53 215 47 48 2 1 2 76 DFFQSRX1 $T=314400 599440 0 0 $X=313970 $Y=599050
X54 85 47 48 2 1 2 89 DFFQSRX1 $T=323360 575920 1 0 $X=322930 $Y=571365
X55 81 47 48 2 1 2 3 DFFQSRX1 $T=349120 568080 1 180 $X=323490 $Y=567690
X56 63 47 48 2 1 2 60 DFFQSRX1 $T=349680 513200 1 180 $X=324050 $Y=512810
X57 78 47 48 2 1 2 4 DFFQSRX1 $T=351360 521040 0 180 $X=325730 $Y=516485
X58 96 47 48 2 1 2 99 DFFQSRX1 $T=341840 536720 1 0 $X=341410 $Y=532165
X59 211 47 48 2 1 2 117 DFFQSRX1 $T=345200 536720 0 0 $X=344770 $Y=536330
X60 125 47 48 2 1 2 118 DFFQSRX1 $T=345200 560240 1 0 $X=344770 $Y=555685
X61 115 47 48 2 1 2 119 DFFQSRX1 $T=345200 560240 0 0 $X=344770 $Y=559850
X62 49 47 48 2 1 2 12 DFFQSRX1 $T=349680 513200 0 0 $X=349250 $Y=512810
X63 95 47 48 2 1 2 10 DFFQSRX1 $T=351360 521040 1 0 $X=350930 $Y=516485
X64 110 47 48 2 1 2 103 DFFQSRX1 $T=386640 568080 1 180 $X=361010 $Y=567690
X65 116 47 48 2 1 2 106 DFFQSRX1 $T=386640 575920 0 180 $X=361010 $Y=571365
X66 121 47 48 2 1 2 123 DFFQSRX1 $T=372080 536720 1 0 $X=371650 $Y=532165
X67 132 47 48 2 1 2 120 DFFQSRX1 $T=397280 536720 1 180 $X=371650 $Y=536330
X68 137 47 48 2 1 2 142 DFFQSRX1 $T=372080 560240 1 0 $X=371650 $Y=555685
X69 122 47 48 2 1 2 126 DFFQSRX1 $T=372080 560240 0 0 $X=371650 $Y=559850
X70 50 47 48 2 1 2 127 DFFQSRX1 $T=376000 513200 0 0 $X=375570 $Y=512810
X71 135 47 48 2 1 2 129 DFFQSRX1 $T=376560 521040 1 0 $X=376130 $Y=516485
X72 145 47 48 2 1 2 138 DFFQSRX1 $T=416880 568080 1 180 $X=391250 $Y=567690
X73 147 47 48 2 1 2 139 DFFQSRX1 $T=416880 575920 0 180 $X=391250 $Y=571365
X74 165 47 48 2 1 2 151 DFFQSRX1 $T=402320 536720 0 0 $X=401890 $Y=536330
X75 146 47 48 2 1 2 152 DFFQSRX1 $T=402320 560240 1 0 $X=401890 $Y=555685
X76 157 47 48 2 1 2 160 DFFQSRX1 $T=403440 536720 1 0 $X=403010 $Y=532165
X77 174 47 48 2 1 2 153 DFFQSRX1 $T=430880 560240 1 180 $X=405250 $Y=559850
X78 167 47 48 2 1 2 173 DFFQSRX1 $T=414640 521040 1 0 $X=414210 $Y=516485
X79 170 47 48 2 1 2 163 DFFQSRX1 $T=442080 568080 1 180 $X=416450 $Y=567690
X80 169 47 48 2 1 2 164 DFFQSRX1 $T=442080 575920 0 180 $X=416450 $Y=571365
X81 51 47 48 2 1 2 21 DFFQSRX1 $T=442640 513200 1 180 $X=417010 $Y=512810
X82 179 47 48 2 1 2 176 DFFQSRX1 $T=458320 536720 1 180 $X=432690 $Y=536330
X83 180 47 48 2 1 2 184 DFFQSRX1 $T=433120 560240 1 0 $X=432690 $Y=555685
X84 194 47 48 2 1 2 182 DFFQSRX1 $T=459440 560240 1 180 $X=433810 $Y=559850
X85 203 47 48 2 1 2 183 DFFQSRX1 $T=461680 536720 0 180 $X=436050 $Y=532165
X86 190 47 48 2 1 2 198 DFFQSRX1 $T=439840 521040 1 0 $X=439410 $Y=516485
X87 186 47 48 2 1 2 191 DFFQSRX1 $T=442080 568080 0 0 $X=441650 $Y=567690
X88 187 47 48 2 1 2 192 DFFQSRX1 $T=442080 575920 1 0 $X=441650 $Y=571365
X89 52 47 48 2 1 2 200 DFFQSRX1 $T=442640 513200 0 0 $X=442210 $Y=512810
X90 199 47 48 2 1 2 204 DFFQSRX1 $T=463360 536720 1 0 $X=462930 $Y=532165
X91 237 47 48 2 1 2 216 DFFQSRX1 $T=491920 536720 1 180 $X=466290 $Y=536330
X92 225 47 48 2 1 2 228 DFFQSRX1 $T=466720 560240 1 0 $X=466290 $Y=555685
X93 227 47 48 2 1 2 234 DFFQSRX1 $T=466720 560240 0 0 $X=466290 $Y=559850
X94 226 47 48 2 1 2 233 DFFQSRX1 $T=474000 568080 0 0 $X=473570 $Y=567690
X95 224 47 48 2 1 2 232 DFFQSRX1 $T=474000 575920 1 0 $X=473570 $Y=571365
X96 241 47 48 2 1 2 221 DFFQSRX1 $T=504800 521040 0 180 $X=479170 $Y=516485
X97 246 47 48 2 1 2 27 DFFQSRX1 $T=508160 513200 1 180 $X=482530 $Y=512810
X98 239 47 48 2 1 2 242 DFFQSRX1 $T=493600 560240 0 0 $X=493170 $Y=559850
X99 254 47 48 2 1 2 253 DFFQSRX1 $T=494720 560240 1 0 $X=494290 $Y=555685
X100 273 47 48 2 1 2 243 DFFQSRX1 $T=522160 536720 0 180 $X=496530 $Y=532165
X101 271 47 48 2 1 2 278 DFFQSRX1 $T=496960 536720 0 0 $X=496530 $Y=536330
X102 255 47 48 2 1 2 258 DFFQSRX1 $T=499200 568080 0 0 $X=498770 $Y=567690
X103 251 47 48 2 1 2 249 DFFQSRX1 $T=499200 575920 1 0 $X=498770 $Y=571365
X104 272 47 48 2 1 2 257 DFFQSRX1 $T=533920 521040 0 180 $X=508290 $Y=516485
X105 54 47 48 2 1 2 31 DFFQSRX1 $T=538400 513200 1 180 $X=512770 $Y=512810
X106 208 47 48 2 1 2 212 DFFQSRX1 $T=524400 536720 1 0 $X=523970 $Y=532165
X107 256 47 48 2 1 2 259 DFFQSRX1 $T=549600 536720 1 180 $X=523970 $Y=536330
X108 268 47 48 2 1 2 263 DFFQSRX1 $T=549600 560240 0 180 $X=523970 $Y=555685
X109 286 47 48 2 1 2 282 DFFQSRX1 $T=552960 560240 1 180 $X=527330 $Y=559850
X110 265 47 48 2 1 2 260 DFFQSRX1 $T=528320 575920 1 0 $X=527890 $Y=571365
X111 280 47 48 2 1 2 266 DFFQSRX1 $T=533920 521040 1 0 $X=533490 $Y=516485
X112 285 47 48 2 1 2 283 DFFQSRX1 $T=534480 568080 0 0 $X=534050 $Y=567690
X113 298 47 48 2 1 2 301 DFFQSRX1 $T=558000 536720 1 0 $X=557570 $Y=532165
X114 292 47 48 2 1 2 295 DFFQSRX1 $T=558000 536720 0 0 $X=557570 $Y=536330
X115 297 47 48 2 1 2 288 DFFQSRX1 $T=583200 560240 0 180 $X=557570 $Y=555685
X116 299 47 48 2 1 2 289 DFFQSRX1 $T=583200 560240 1 180 $X=557570 $Y=559850
X117 290 47 48 2 1 2 291 DFFQSRX1 $T=558560 575920 1 0 $X=558130 $Y=571365
X118 293 47 48 2 1 2 296 DFFQSRX1 $T=559680 568080 0 0 $X=559250 $Y=567690
X119 1 47 48 2 1 2 37 DFFQSRX1 $T=560240 513200 0 0 $X=559810 $Y=512810
X120 1 47 48 2 1 2 38 DFFQSRX1 $T=561360 521040 1 0 $X=560930 $Y=516485
X121 302 47 48 2 1 2 300 DFFQSRX1 $T=584880 536720 0 0 $X=584450 $Y=536330
X122 307 47 48 2 1 2 312 DFFQSRX1 $T=586000 560240 1 0 $X=585570 $Y=555685
X123 303 47 48 2 1 2 310 DFFQSRX1 $T=586560 536720 1 0 $X=586130 $Y=532165
X124 306 47 48 2 1 2 311 DFFQSRX1 $T=586560 560240 0 0 $X=586130 $Y=559850
X125 308 47 48 2 1 2 315 DFFQSRX1 $T=588800 568080 0 0 $X=588370 $Y=567690
X126 309 47 48 2 1 2 294 DFFQSRX1 $T=588800 575920 1 0 $X=588370 $Y=571365
X127 320 47 48 2 1 2 316 DFFQSRX1 $T=593840 521040 1 0 $X=593410 $Y=516485
X128 322 47 48 2 1 2 314 DFFQSRX1 $T=624080 513200 1 180 $X=598450 $Y=512810
X129 328 47 48 2 1 2 323 DFFQSRX1 $T=640880 560240 0 180 $X=615250 $Y=555685
X130 327 47 48 2 1 2 329 DFFQSRX1 $T=619600 544560 1 0 $X=619170 $Y=540005
X131 321 47 48 2 1 2 324 DFFQSRX1 $T=619600 575920 1 0 $X=619170 $Y=571365
X132 331 47 48 2 1 2 325 DFFQSRX1 $T=619600 583760 1 0 $X=619170 $Y=579205
X133 318 47 48 2 1 2 304 DFFQSRX1 $T=619600 583760 0 0 $X=619170 $Y=583370
X134 326 47 48 2 1 2 317 DFFQSRX1 $T=619600 599440 1 0 $X=619170 $Y=594885
X135 287 47 48 2 1 2 284 DFFQSRX1 $T=619600 599440 0 0 $X=619170 $Y=599050
X136 349 47 48 2 1 2 330 DFFQSRX1 $T=624640 591600 0 0 $X=624210 $Y=591210
X137 338 47 48 2 1 2 339 DFFQSRX1 $T=628000 552400 0 0 $X=627570 $Y=552010
X138 342 47 48 2 1 2 45 DFFQSRX1 $T=654320 505360 1 180 $X=628690 $Y=504970
X139 343 47 48 2 1 2 332 DFFQSRX1 $T=654320 521040 0 180 $X=628690 $Y=516485
X140 344 47 48 2 1 2 333 DFFQSRX1 $T=654320 528880 0 180 $X=628690 $Y=524325
X141 345 47 48 2 1 2 334 DFFQSRX1 $T=654320 536720 0 180 $X=628690 $Y=532165
X142 346 47 48 2 1 2 335 DFFQSRX1 $T=654320 544560 1 180 $X=628690 $Y=544170
X143 340 47 48 2 1 2 341 DFFQSRX1 $T=629120 575920 0 0 $X=628690 $Y=575530
X144 348 47 48 2 1 2 336 DFFQSRX1 $T=654320 591600 0 180 $X=628690 $Y=587045
X145 347 47 48 2 1 2 337 DFFQSRX1 $T=654880 568080 0 180 $X=629250 $Y=563525
X277 62 3 1 2 61 NAND2X1 $T=335680 568080 0 180 $X=332450 $Y=563525
X278 67 71 1 2 70 NAND2X1 $T=335680 591600 1 0 $X=335250 $Y=587045
X279 5 75 1 2 77 NAND2X1 $T=337920 575920 0 0 $X=337490 $Y=575530
X280 80 75 1 2 67 NAND2X1 $T=343520 591600 0 180 $X=340290 $Y=587045
X281 7 61 1 2 81 NAND2X1 $T=345200 568080 0 180 $X=341970 $Y=563525
X282 89 9 1 2 88 NAND2X1 $T=348000 568080 1 0 $X=347570 $Y=563525
X283 91 90 1 2 80 NAND2X1 $T=350800 583760 1 180 $X=347570 $Y=583370
X284 93 94 1 2 62 NAND2X1 $T=354720 575920 0 180 $X=351490 $Y=571365
X285 103 94 1 2 100 NAND2X1 $T=358640 575920 0 0 $X=358210 $Y=575530
X286 112 94 1 2 111 NAND2X1 $T=366480 568080 0 180 $X=363250 $Y=563525
X287 114 94 1 2 113 NAND2X1 $T=367040 583760 0 180 $X=363810 $Y=579205
X288 103 108 1 2 114 NAND2X1 $T=367040 583760 1 180 $X=363810 $Y=583370
X289 109 106 1 2 87 NAND2X1 $T=364800 591600 1 0 $X=364370 $Y=587045
X290 103 9 1 2 112 NAND2X1 $T=366480 568080 1 0 $X=366050 $Y=563525
X291 13 120 1 2 124 NAND2X1 $T=379360 544560 0 180 $X=376130 $Y=540005
X292 13 127 1 2 14 NAND2X1 $T=379920 513200 1 0 $X=379490 $Y=508645
X293 13 129 1 2 128 NAND2X1 $T=380480 528880 0 0 $X=380050 $Y=528490
X294 16 129 1 2 15 NAND2X1 $T=386080 521040 1 180 $X=382850 $Y=520650
X295 16 127 1 2 131 NAND2X1 $T=386080 528880 1 180 $X=382850 $Y=528490
X296 16 120 1 2 133 NAND2X1 $T=390560 544560 0 180 $X=387330 $Y=540005
X297 17 123 1 2 134 NAND2X1 $T=394480 528880 1 180 $X=391250 $Y=528490
X298 13 142 1 2 141 NAND2X1 $T=391680 544560 1 0 $X=391250 $Y=540005
X299 16 56 1 2 18 NAND2X1 $T=394480 521040 0 0 $X=394050 $Y=520650
X300 17 118 1 2 140 NAND2X1 $T=400080 544560 1 180 $X=396850 $Y=544170
X301 16 142 1 2 136 NAND2X1 $T=400640 536720 1 180 $X=397410 $Y=536330
X302 17 126 1 2 130 NAND2X1 $T=397840 544560 1 0 $X=397410 $Y=540005
X303 13 56 1 2 144 NAND2X1 $T=401760 521040 1 180 $X=398530 $Y=520650
X304 16 151 1 2 150 NAND2X1 $T=403440 544560 1 0 $X=403010 $Y=540005
X305 17 152 1 2 154 NAND2X1 $T=406800 544560 1 0 $X=406370 $Y=540005
X306 17 72 1 2 148 NAND2X1 $T=408480 521040 1 0 $X=408050 $Y=516485
X307 17 138 1 2 156 NAND2X1 $T=411840 544560 1 180 $X=408610 $Y=544170
X308 16 20 1 2 155 NAND2X1 $T=411840 521040 1 0 $X=411410 $Y=516485
X309 13 151 1 2 159 NAND2X1 $T=414640 544560 1 180 $X=411410 $Y=544170
X310 13 20 1 2 19 NAND2X1 $T=412400 505360 0 0 $X=411970 $Y=504970
X311 13 160 1 2 158 NAND2X1 $T=412400 528880 0 0 $X=411970 $Y=528490
X312 17 139 1 2 162 NAND2X1 $T=414640 544560 0 0 $X=414210 $Y=544170
X313 16 160 1 2 161 NAND2X1 $T=415200 528880 0 0 $X=414770 $Y=528490
X314 17 163 1 2 168 NAND2X1 $T=420240 544560 0 0 $X=419810 $Y=544170
X315 13 153 1 2 172 NAND2X1 $T=425280 552400 0 180 $X=422050 $Y=547845
X316 16 153 1 2 166 NAND2X1 $T=426960 544560 0 180 $X=423730 $Y=540005
X317 16 173 1 2 22 NAND2X1 $T=424720 521040 0 0 $X=424290 $Y=520650
X318 16 176 1 2 175 NAND2X1 $T=426960 544560 1 0 $X=426530 $Y=540005
X319 13 173 1 2 171 NAND2X1 $T=428640 536720 1 0 $X=428210 $Y=532165
X320 17 164 1 2 177 NAND2X1 $T=432000 552400 0 180 $X=428770 $Y=547845
X321 16 21 1 2 178 NAND2X1 $T=433680 521040 1 180 $X=430450 $Y=520650
X322 13 176 1 2 181 NAND2X1 $T=435360 544560 0 180 $X=432130 $Y=540005
X323 16 182 1 2 185 NAND2X1 $T=442080 544560 1 0 $X=441650 $Y=540005
X324 17 184 1 2 188 NAND2X1 $T=444320 544560 0 0 $X=443890 $Y=544170
X325 13 182 1 2 189 NAND2X1 $T=449920 544560 0 180 $X=446690 $Y=540005
X326 16 198 1 2 23 NAND2X1 $T=449920 528880 1 0 $X=449490 $Y=524325
X327 13 183 1 2 197 NAND2X1 $T=450480 544560 1 0 $X=450050 $Y=540005
X328 17 192 1 2 193 NAND2X1 $T=453280 552400 0 180 $X=450050 $Y=547845
X329 16 183 1 2 196 NAND2X1 $T=454960 544560 1 180 $X=451730 $Y=544170
X330 13 198 1 2 195 NAND2X1 $T=452720 528880 1 0 $X=452290 $Y=524325
X331 13 200 1 2 24 NAND2X1 $T=454400 505360 0 0 $X=453970 $Y=504970
X332 16 200 1 2 202 NAND2X1 $T=456080 528880 1 0 $X=455650 $Y=524325
X333 17 191 1 2 201 NAND2X1 $T=456640 544560 0 0 $X=456210 $Y=544170
X334 16 58 1 2 206 NAND2X1 $T=459440 544560 0 0 $X=459010 $Y=544170
X335 16 212 1 2 25 NAND2X1 $T=461680 528880 1 0 $X=461250 $Y=524325
X336 13 212 1 2 210 NAND2X1 $T=462800 536720 0 0 $X=462370 $Y=536330
X337 13 117 1 2 214 NAND2X1 $T=463360 544560 0 0 $X=462930 $Y=544170
X338 16 117 1 2 205 NAND2X1 $T=465600 544560 1 0 $X=465170 $Y=540005
X339 17 74 1 2 213 NAND2X1 $T=468960 544560 1 180 $X=465730 $Y=544170
X340 17 204 1 2 207 NAND2X1 $T=468960 544560 1 0 $X=468530 $Y=540005
X341 17 76 1 2 217 NAND2X1 $T=468960 544560 0 0 $X=468530 $Y=544170
X342 13 58 1 2 218 NAND2X1 $T=474560 544560 0 180 $X=471330 $Y=540005
X343 16 26 1 2 219 NAND2X1 $T=476240 521040 1 180 $X=473010 $Y=520650
X344 13 216 1 2 223 NAND2X1 $T=481840 528880 0 0 $X=481410 $Y=528490
X345 13 228 1 2 222 NAND2X1 $T=481840 544560 1 0 $X=481410 $Y=540005
X346 13 221 1 2 230 NAND2X1 $T=483520 521040 0 0 $X=483090 $Y=520650
X347 16 216 1 2 231 NAND2X1 $T=487440 544560 0 180 $X=484210 $Y=540005
X348 16 221 1 2 28 NAND2X1 $T=489120 521040 1 180 $X=485890 $Y=520650
X349 17 234 1 2 229 NAND2X1 $T=490800 544560 1 180 $X=487570 $Y=544170
X350 16 228 1 2 235 NAND2X1 $T=491360 536720 0 180 $X=488130 $Y=532165
X351 16 29 1 2 238 NAND2X1 $T=490240 521040 0 0 $X=489810 $Y=520650
X352 17 233 1 2 236 NAND2X1 $T=493600 544560 1 180 $X=490370 $Y=544170
X353 17 232 1 2 240 NAND2X1 $T=492480 544560 1 0 $X=492050 $Y=540005
X354 13 29 1 2 30 NAND2X1 $T=496960 513200 0 180 $X=493730 $Y=508645
X355 17 242 1 2 244 NAND2X1 $T=498640 544560 0 180 $X=495410 $Y=540005
X356 17 249 1 2 247 NAND2X1 $T=497520 544560 0 0 $X=497090 $Y=544170
X357 13 27 1 2 248 NAND2X1 $T=498080 513200 1 0 $X=497650 $Y=508645
X358 13 253 1 2 252 NAND2X1 $T=501440 544560 1 0 $X=501010 $Y=540005
X359 16 243 1 2 250 NAND2X1 $T=503120 528880 0 0 $X=502690 $Y=528490
X360 16 253 1 2 245 NAND2X1 $T=505920 528880 0 0 $X=505490 $Y=528490
X361 17 259 1 2 261 NAND2X1 $T=511520 521040 0 0 $X=511090 $Y=520650
X362 17 263 1 2 262 NAND2X1 $T=512080 528880 0 0 $X=511650 $Y=528490
X363 13 243 1 2 264 NAND2X1 $T=515440 544560 0 180 $X=512210 $Y=540005
X364 16 266 1 2 32 NAND2X1 $T=514880 513200 1 0 $X=514450 $Y=508645
X365 17 260 1 2 267 NAND2X1 $T=518240 544560 0 180 $X=515010 $Y=540005
X366 16 257 1 2 269 NAND2X1 $T=517680 521040 0 0 $X=517250 $Y=520650
X367 16 33 1 2 270 NAND2X1 $T=522160 513200 0 180 $X=518930 $Y=508645
X368 16 278 1 2 276 NAND2X1 $T=520480 521040 0 0 $X=520050 $Y=520650
X369 16 31 1 2 279 NAND2X1 $T=522160 513200 1 0 $X=521730 $Y=508645
X370 13 278 1 2 275 NAND2X1 $T=525520 544560 0 180 $X=522290 $Y=540005
X371 13 257 1 2 277 NAND2X1 $T=528320 528880 0 180 $X=525090 $Y=524325
X372 17 258 1 2 274 NAND2X1 $T=528320 544560 0 180 $X=525090 $Y=540005
X373 13 266 1 2 281 NAND2X1 $T=526080 513200 1 0 $X=525650 $Y=508645
X374 35 305 1 2 313 NAND2X1 $T=600000 528880 0 180 $X=596770 $Y=524325
X375 314 316 1 2 43 NAND2X1 $T=598320 513200 1 0 $X=597890 $Y=508645
X376 44 316 1 2 319 NAND2X1 $T=606160 513200 0 180 $X=602930 $Y=508645
X377 319 313 1 2 320 NAND2X1 $T=606160 521040 1 180 $X=602930 $Y=520650
X460 87 103 1 2 101 AND2X1 $T=362000 583760 1 180 $X=358210 $Y=583370
X461 119 11 1 2 109 AND2X1 $T=371520 583760 1 0 $X=371090 $Y=579205
X462 60 5 6 1 2 63 MUX2X1 $T=341280 505360 1 180 $X=335250 $Y=504970
X463 73 5 60 1 2 64 MUX2X1 $T=341280 528880 1 180 $X=335250 $Y=528490
X464 73 7 68 1 2 65 MUX2X1 $T=341280 544560 1 180 $X=335250 $Y=544170
X465 57 5 73 1 2 79 MUX2X1 $T=335680 552400 1 0 $X=335250 $Y=547845
X466 57 7 69 1 2 66 MUX2X1 $T=341280 568080 0 180 $X=335250 $Y=563525
X467 4 5 57 1 2 78 MUX2X1 $T=345200 528880 0 180 $X=339170 $Y=524325
X468 97 59 91 1 2 102 MUX2X1 $T=350800 591600 1 0 $X=350370 $Y=587045
X469 60 7 10 1 2 95 MUX2X1 $T=357520 513200 0 180 $X=351490 $Y=508645
X470 4 7 99 1 2 96 MUX2X1 $T=357520 521040 1 180 $X=351490 $Y=520650
X471 5 119 111 1 2 115 MUX2X1 $T=373760 575920 1 180 $X=367730 $Y=575530
X472 107 106 113 1 2 116 MUX2X1 $T=374880 591600 0 180 $X=368850 $Y=587045
X473 123 3 99 1 2 121 MUX2X1 $T=378800 528880 1 180 $X=372770 $Y=528490
X474 126 3 68 1 2 122 MUX2X1 $T=381600 552400 1 180 $X=375570 $Y=552010
X475 118 3 69 1 2 125 MUX2X1 $T=384400 568080 0 180 $X=378370 $Y=563525
X476 72 3 123 1 2 143 MUX2X1 $T=402320 528880 1 180 $X=396290 $Y=528490
X477 138 3 126 1 2 145 MUX2X1 $T=405680 560240 1 180 $X=399650 $Y=559850
X478 152 3 72 1 2 146 MUX2X1 $T=407360 544560 1 180 $X=401330 $Y=544170
X479 139 3 118 1 2 147 MUX2X1 $T=408480 575920 1 180 $X=402450 $Y=575530
X480 164 3 138 1 2 169 MUX2X1 $T=427520 568080 0 180 $X=421490 $Y=563525
X481 163 3 139 1 2 170 MUX2X1 $T=427520 583760 0 180 $X=421490 $Y=579205
X482 184 3 152 1 2 180 MUX2X1 $T=438160 552400 0 180 $X=432130 $Y=547845
X483 191 3 164 1 2 186 MUX2X1 $T=448800 575920 1 180 $X=442770 $Y=575530
X484 192 3 163 1 2 187 MUX2X1 $T=448800 583760 1 180 $X=442770 $Y=583370
X485 204 3 184 1 2 199 MUX2X1 $T=459440 552400 1 180 $X=453410 $Y=552010
X486 74 3 192 1 2 209 MUX2X1 $T=467280 583760 0 180 $X=461250 $Y=579205
X487 76 3 191 1 2 215 MUX2X1 $T=471200 575920 1 180 $X=465170 $Y=575530
X488 232 3 204 1 2 224 MUX2X1 $T=488560 568080 0 180 $X=482530 $Y=563525
X489 233 3 76 1 2 226 MUX2X1 $T=489120 575920 1 180 $X=483090 $Y=575530
X490 234 3 74 1 2 227 MUX2X1 $T=489120 583760 1 180 $X=483090 $Y=583370
X491 242 3 232 1 2 239 MUX2X1 $T=496960 552400 1 180 $X=490930 $Y=552010
X492 249 3 234 1 2 251 MUX2X1 $T=508160 575920 1 180 $X=502130 $Y=575530
X493 258 3 233 1 2 255 MUX2X1 $T=510400 568080 0 180 $X=504370 $Y=563525
X494 259 3 242 1 2 256 MUX2X1 $T=512080 544560 0 180 $X=506050 $Y=540005
X495 260 3 249 1 2 265 MUX2X1 $T=510400 575920 0 0 $X=509970 $Y=575530
X496 263 3 258 1 2 268 MUX2X1 $T=512640 568080 1 0 $X=512210 $Y=563525
X497 283 35 282 1 2 285 MUX2X1 $T=545120 575920 0 0 $X=544690 $Y=575530
X498 282 35 284 1 2 286 MUX2X1 $T=545120 591600 1 0 $X=544690 $Y=587045
X499 36 35 283 1 2 34 MUX2X1 $T=551280 568080 0 180 $X=545250 $Y=563525
X500 284 35 288 1 2 287 MUX2X1 $T=556320 591600 0 180 $X=550290 $Y=587045
X501 291 35 36 1 2 290 MUX2X1 $T=568640 568080 0 180 $X=562610 $Y=563525
X502 295 35 289 1 2 292 MUX2X1 $T=574240 552400 1 180 $X=568210 $Y=552010
X503 288 35 296 1 2 297 MUX2X1 $T=569200 591600 1 0 $X=568770 $Y=587045
X504 289 35 291 1 2 299 MUX2X1 $T=569760 568080 1 0 $X=569330 $Y=563525
X505 296 35 294 1 2 293 MUX2X1 $T=575360 583760 0 180 $X=569330 $Y=579205
X506 301 35 300 1 2 298 MUX2X1 $T=580400 528880 1 180 $X=574370 $Y=528490
X507 300 35 295 1 2 302 MUX2X1 $T=574800 552400 0 0 $X=574370 $Y=552010
X508 294 35 304 1 2 309 MUX2X1 $T=591040 583760 1 0 $X=590610 $Y=579205
X509 310 35 301 1 2 303 MUX2X1 $T=599440 528880 1 180 $X=593410 $Y=528490
X510 311 35 310 1 2 306 MUX2X1 $T=601680 544560 0 180 $X=595650 $Y=540005
X511 312 35 311 1 2 307 MUX2X1 $T=601680 544560 1 180 $X=595650 $Y=544170
X512 315 35 312 1 2 308 MUX2X1 $T=601680 568080 0 180 $X=595650 $Y=563525
X513 304 35 317 1 2 318 MUX2X1 $T=598880 583760 1 0 $X=598450 $Y=579205
X514 35 314 44 1 2 322 MUX2X1 $T=608400 513200 1 0 $X=607970 $Y=508645
X515 324 35 315 1 2 321 MUX2X1 $T=618480 568080 0 180 $X=612450 $Y=563525
X516 317 35 325 1 2 326 MUX2X1 $T=612880 591600 1 0 $X=612450 $Y=587045
X517 323 35 324 1 2 328 MUX2X1 $T=618480 568080 1 0 $X=618050 $Y=563525
X518 329 35 323 1 2 327 MUX2X1 $T=625760 552400 1 180 $X=619730 $Y=552010
X519 325 35 330 1 2 331 MUX2X1 $T=620720 591600 1 0 $X=620290 $Y=587045
X520 339 35 329 1 2 338 MUX2X1 $T=636960 552400 0 180 $X=630930 $Y=547845
X521 45 35 332 1 2 342 MUX2X1 $T=639200 513200 1 0 $X=638770 $Y=508645
X522 332 35 333 1 2 343 MUX2X1 $T=639200 521040 0 0 $X=638770 $Y=520650
X523 333 35 334 1 2 344 MUX2X1 $T=639200 528880 0 0 $X=638770 $Y=528490
X524 334 35 335 1 2 345 MUX2X1 $T=639200 536720 0 0 $X=638770 $Y=536330
X525 335 35 339 1 2 346 MUX2X1 $T=639200 552400 1 0 $X=638770 $Y=547845
X526 341 35 337 1 2 340 MUX2X1 $T=644800 568080 1 180 $X=638770 $Y=567690
X527 337 35 46 1 2 347 MUX2X1 $T=644800 575920 1 0 $X=644370 $Y=571365
X528 336 35 341 1 2 348 MUX2X1 $T=644800 583760 1 0 $X=644370 $Y=579205
X529 330 35 336 1 2 349 MUX2X1 $T=644800 583760 0 0 $X=644370 $Y=583370
X530 83 9 1 2 98 NOR2X1 $T=351360 568080 1 0 $X=350930 $Y=563525
X531 89 101 1 2 91 NOR2X1 $T=354160 583760 1 0 $X=353730 $Y=579205
X532 9 100 1 2 5 NOR2X1 $T=360320 568080 1 0 $X=359890 $Y=563525
X533 108 100 1 2 107 NOR2X1 $T=363680 591600 1 180 $X=360450 $Y=591210
X534 41 43 1 2 42 NOR2X1 $T=596080 505360 0 0 $X=595650 $Y=504970
X535 75 1 2 82 INVX2 $T=342960 583760 0 0 $X=342530 $Y=583370
X536 8 1 2 83 INVX2 $T=343520 536720 0 0 $X=343090 $Y=536330
X537 100 1 2 92 INVX2 $T=353040 591600 0 0 $X=352610 $Y=591210
X538 103 1 2 93 INVX2 $T=356960 575920 0 180 $X=354850 $Y=571365
X539 89 1 2 94 INVX2 $T=356960 575920 1 180 $X=354850 $Y=575530
X540 109 1 2 108 INVX2 $T=364240 583760 1 180 $X=362130 $Y=583370
X541 11 1 2 9 INVX2 $T=451600 552400 1 180 $X=449490 $Y=552010
X542 40 1 2 39 INVX2 $T=592160 505360 1 180 $X=590050 $Y=504970
X729 77 86 88 1 2 85 NAND3X1 $T=343520 575920 0 0 $X=343090 $Y=575530
X730 92 59 82 1 2 84 NAND3X1 $T=350800 591600 0 180 $X=346450 $Y=587045
X731 93 94 83 1 2 86 NAND3X1 $T=354160 575920 1 180 $X=349810 $Y=575530
X732 103 89 98 1 2 7 NAND3X1 $T=358080 568080 0 180 $X=353730 $Y=563525
X733 93 89 11 1 2 105 NAND3X1 $T=356960 575920 1 0 $X=356530 $Y=571365
X734 112 100 105 1 2 110 NAND3X1 $T=366480 575920 1 180 $X=362130 $Y=575530
X735 124 130 131 1 2 132 NAND3X1 $T=381600 544560 1 0 $X=381170 $Y=540005
X736 128 134 136 1 2 135 NAND3X1 $T=387760 528880 0 0 $X=387330 $Y=528490
X737 141 140 133 1 2 137 NAND3X1 $T=394480 544560 1 180 $X=390130 $Y=544170
X738 144 148 150 1 2 149 NAND3X1 $T=401760 521040 1 0 $X=401330 $Y=516485
X739 158 156 155 1 2 157 NAND3X1 $T=413520 544560 0 180 $X=409170 $Y=540005
X740 159 162 161 1 2 165 NAND3X1 $T=414640 544560 1 0 $X=414210 $Y=540005
X741 171 154 166 1 2 167 NAND3X1 $T=424160 544560 0 180 $X=419810 $Y=540005
X742 172 168 175 1 2 174 NAND3X1 $T=425280 552400 1 0 $X=424850 $Y=547845
X743 181 177 178 1 2 179 NAND3X1 $T=435360 536720 0 180 $X=431010 $Y=532165
X744 189 193 196 1 2 194 NAND3X1 $T=445440 552400 1 0 $X=445010 $Y=547845
X745 195 188 185 1 2 190 NAND3X1 $T=449920 528880 1 180 $X=445570 $Y=528490
X746 197 201 202 1 2 203 NAND3X1 $T=454960 544560 1 0 $X=454530 $Y=540005
X747 210 207 205 1 2 208 NAND3X1 $T=463920 544560 0 180 $X=459570 $Y=540005
X748 214 213 206 1 2 211 NAND3X1 $T=466160 552400 1 180 $X=461810 $Y=552010
X749 218 217 219 1 2 220 NAND3X1 $T=471760 544560 0 0 $X=471330 $Y=544170
X750 222 229 231 1 2 225 NAND3X1 $T=481840 544560 0 0 $X=481410 $Y=544170
X751 223 236 238 1 2 237 NAND3X1 $T=488000 544560 1 0 $X=487570 $Y=540005
X752 230 240 235 1 2 241 NAND3X1 $T=490800 528880 0 0 $X=490370 $Y=528490
X753 248 244 245 1 2 246 NAND3X1 $T=501440 528880 1 180 $X=497090 $Y=528490
X754 252 247 250 1 2 254 NAND3X1 $T=506480 544560 1 180 $X=502130 $Y=544170
X755 275 267 269 1 2 271 NAND3X1 $T=522160 544560 1 180 $X=517810 $Y=544170
X756 277 262 270 1 2 272 NAND3X1 $T=522720 528880 0 180 $X=518370 $Y=524325
X757 264 274 279 1 2 273 NAND3X1 $T=518800 544560 1 0 $X=518370 $Y=540005
X758 281 261 276 1 2 280 NAND3X1 $T=529440 521040 1 180 $X=525090 $Y=520650
X776 87 84 1 2 71 OR2X1 $T=346880 591600 0 180 $X=343090 $Y=587045
X777 93 59 1 2 90 OR2X1 $T=351920 575920 0 180 $X=348130 $Y=571365
X778 100 87 1 2 97 OR2X1 $T=360880 591600 0 180 $X=357090 $Y=587045
X779 316 314 2 1 305 XOR2X1 $T=601680 521040 1 180 $X=595090 $Y=520650
X780 102 1 2 104 INVX1 $T=356960 591600 0 0 $X=356530 $Y=591210
.ENDS
***************************************
.SUBCKT ICV_35
** N=4 EP=0 IP=1 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=4 EP=0 IP=72 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4
** N=6 EP=4 IP=6 FDC=96
X0 1 4 2 3 pad_in $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4
** N=6 EP=4 IP=6 FDC=96
X0 1 4 2 3 pad_in $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4
** N=6 EP=4 IP=6 FDC=96
X0 1 4 2 3 pad_in $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_2 VSS VDD
** N=46 EP=2 IP=1 FDC=1
D0 VSS VDD ndio_m AREA=9e-10 PJ=0.00012 $X=10780 $Y=193610 $D=30
.ENDS
***************************************
.SUBCKT ICV_31
** N=5 EP=0 IP=44 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=4 EP=0 IP=72 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28
** N=4 EP=0 IP=72 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=4 EP=0 IP=72 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=4 EP=0 IP=40 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4
** N=6 EP=4 IP=6 FDC=96
X0 2 3 4 1 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4
** N=6 EP=4 IP=6 FDC=96
X0 1 4 2 3 pad_in $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT bridge_soc_top VSS VDD Bridge_Serial_out Serial_in clock T_byte R_byte reset Bridge_Can_out Can_rx
** N=153 EP=10 IP=459 FDC=17522
X3 VSS VDD 3 Bridge_Serial_out ICV_12 $T=0 413840 0 270 $X=0 $Y=322940
X6 VSS VDD 4 Serial_in ICV_8 $T=0 594480 0 270 $X=0 $Y=503580
X22 VSS VDD ICV_1 $T=291700 0 0 0 $X=290800 $Y=0
X23 VSS VDD clock ICV_4 $T=381700 918320 0 180 $X=290800 $Y=684220
X26 VSS VDD 12 14 7 10 11 16 17 78 18 20 19 21 22 23 24 26 25 27
+ 29 6 30 77 13 15 8 28
+ ICV_52 $T=0 0 0 0 $X=292300 $Y=264600
X27 61 VSS VDD 3 80 31 51 79 100 62 102 8 9 7 32 10 12 11 13 103
+ 33 14 34 15 105 21 17 35 82 16 106 107 54 18 88 19 108 20 89 90
+ 109 37 83 112 93 111 110 115 38 91 113 92 39 118 116 40 94 117 95 119
+ 120 121 22 42 122 123 43 24 25 23 96 5 26 29 27 98 124 28 125 99
+ 85 77 30 86 101 87 81 104 78 36 114 41 97 84
+ ICV_51 $T=0 0 0 0 $X=292300 $Y=324400
X28 VSS VDD 44 31 32 4 45 126 79 127 47 48 100 51 46 86 101 62 80 103
+ 128 87 129 34 61 33 130 102 131 104 105 81 82 49 35 52 132 50 54 106
+ 53 88 36 107 89 90 133 91 109 134 55 83 37 56 135 57 92 114 113 58
+ 39 136 115 38 59 93 60 116 118 117 94 63 41 64 40 137 119 120 95 65
+ 66 121 122 68 67 75 138 42 123 125 69 70 96 71 140 73 97 72 43 84
+ 124 98 99 74 77 30 110 108 111 112 139
+ ICV_47 $T=0 0 0 0 $X=292300 $Y=430200
X29 VSS VDD 79 47 45 44 126 4 138 46 75 127 51 129 130 62 61 131 49 50
+ 52 132 133 55 135 57 60 136 58 59 65 63 137 139 125 66 67 68 71 73
+ 70 72 140 69 74 76 77 30 48 128 53 134 64
+ ICV_45 $T=0 0 0 0 $X=292300 $Y=504970
X33 VSS VDD 5 T_byte ICV_14 $T=440200 0 0 0 $X=439300 $Y=0
X34 VSS VDD 75 R_byte ICV_3 $T=530200 918320 0 180 $X=439300 $Y=684220
X35 VSS VDD 6 reset ICV_13 $T=588700 0 0 0 $X=587800 $Y=0
X36 VSS VDD ICV_2 $T=678700 918320 0 180 $X=587800 $Y=684220
X46 VSS VDD 85 Bridge_Can_out ICV_11 $T=970400 323840 0 90 $X=736300 $Y=322940
X48 VSS VDD 76 Can_rx ICV_7 $T=970400 504480 0 90 $X=736300 $Y=503580
.ENDS
***************************************
