/research/ece/lnis-teaching/Designkits/tsmc180nm/full_custom_lib/lef/tech.lef